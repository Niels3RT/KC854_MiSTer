library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_m026 is
    generic(
        ADDR_WIDTH   : integer := 13
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom_m026;

architecture rtl of rom_m026 is
    type rom8192x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom8192x8 := (
         x"7f",  x"7f",  x"46",  x"4f",  x"52",  x"54",  x"48",  x"01", -- 0000
         x"c3",  x"cc",  x"d8",  x"7f",  x"7f",  x"52",  x"45",  x"46", -- 0008
         x"4f",  x"52",  x"54",  x"48",  x"00",  x"c3",  x"b6",  x"d8", -- 0010
         x"00",  x"c3",  x"cc",  x"d8",  x"00",  x"c3",  x"b6",  x"d8", -- 0018
         x"03",  x"00",  x"01",  x"00",  x"10",  x"c9",  x"08",  x"00", -- 0020
         x"00",  x"02",  x"e0",  x"00",  x"7e",  x"01",  x"e0",  x"00", -- 0028
         x"1f",  x"00",  x"00",  x"00",  x"8d",  x"02",  x"8d",  x"02", -- 0030
         x"8b",  x"02",  x"f0",  x"2f",  x"00",  x"40",  x"00",  x"04", -- 0038
         x"00",  x"00",  x"84",  x"43",  x"41",  x"4f",  x"d3",  x"cd", -- 0040
         x"df",  x"4b",  x"c0",  x"e1",  x"d1",  x"c5",  x"cd",  x"0c", -- 0048
         x"f0",  x"c1",  x"c3",  x"1b",  x"c9",  x"86",  x"4e",  x"4f", -- 0050
         x"52",  x"4d",  x"49",  x"ce",  x"42",  x"c0",  x"d8",  x"cd", -- 0058
         x"2c",  x"c9",  x"48",  x"02",  x"64",  x"cd",  x"2c",  x"c9", -- 0060
         x"bb",  x"b7",  x"0b",  x"c1",  x"2c",  x"c9",  x"04",  x"00", -- 0068
         x"2b",  x"cf",  x"d6",  x"cf",  x"a4",  x"cd",  x"18",  x"cc", -- 0070
         x"87",  x"4e",  x"4f",  x"52",  x"4d",  x"4f",  x"55",  x"d4", -- 0078
         x"55",  x"c0",  x"d8",  x"cd",  x"2c",  x"c9",  x"20",  x"00", -- 0080
         x"56",  x"ce",  x"49",  x"c0",  x"56",  x"ce",  x"2b",  x"cf", -- 0088
         x"a4",  x"cd",  x"18",  x"cc",  x"85",  x"53",  x"45",  x"54", -- 0090
         x"49",  x"ce",  x"78",  x"c0",  x"d8",  x"cd",  x"2b",  x"cf", -- 0098
         x"d6",  x"cf",  x"2c",  x"c9",  x"1f",  x"00",  x"fa",  x"cc", -- 00A0
         x"49",  x"c0",  x"a4",  x"cd",  x"18",  x"cc",  x"86",  x"53", -- 00A8
         x"45",  x"54",  x"4f",  x"55",  x"d4",  x"94",  x"c0",  x"d8", -- 00B0
         x"cd",  x"2b",  x"cf",  x"2c",  x"c9",  x"1e",  x"00",  x"fa", -- 00B8
         x"cc",  x"49",  x"c0",  x"a4",  x"cd",  x"18",  x"cc",  x"83", -- 00C0
         x"49",  x"43",  x"c0",  x"ae",  x"c0",  x"cf",  x"c0",  x"e1", -- 00C8
         x"1e",  x"29",  x"cd",  x"0c",  x"f0",  x"6f",  x"26",  x"00", -- 00D0
         x"c3",  x"1a",  x"c9",  x"82",  x"49",  x"c0",  x"c7",  x"c0", -- 00D8
         x"e2",  x"c0",  x"e1",  x"1e",  x"29",  x"cd",  x"0c",  x"f0", -- 00E0
         x"57",  x"23",  x"cd",  x"0c",  x"f0",  x"5a",  x"57",  x"d5", -- 00E8
         x"c3",  x"1b",  x"c9",  x"83",  x"49",  x"43",  x"a1",  x"db", -- 00F0
         x"c0",  x"fb",  x"c0",  x"e1",  x"d1",  x"7b",  x"1e",  x"28", -- 00F8
         x"cd",  x"0c",  x"f0",  x"c3",  x"1b",  x"c9",  x"82",  x"49", -- 0100
         x"a1",  x"f3",  x"c0",  x"0d",  x"c1",  x"e1",  x"d1",  x"7b", -- 0108
         x"1e",  x"28",  x"cd",  x"0c",  x"f0",  x"7a",  x"23",  x"cd", -- 0110
         x"0c",  x"f0",  x"c3",  x"1b",  x"c9",  x"83",  x"42",  x"59", -- 0118
         x"c5",  x"06",  x"c1",  x"d8",  x"cd",  x"5e",  x"c0",  x"82", -- 0120
         x"c0",  x"fa",  x"ca",  x"2c",  x"c9",  x"12",  x"00",  x"56", -- 0128
         x"ce",  x"49",  x"c0",  x"18",  x"cc",  x"86",  x"53",  x"57", -- 0130
         x"49",  x"54",  x"43",  x"c8",  x"1d",  x"c1",  x"40",  x"c1", -- 0138
         x"e1",  x"d1",  x"53",  x"1e",  x"26",  x"3e",  x"02",  x"cd", -- 0140
         x"0c",  x"f0",  x"c3",  x"1b",  x"c9",  x"85",  x"4d",  x"4f", -- 0148
         x"44",  x"55",  x"cc",  x"35",  x"c1",  x"57",  x"c1",  x"e1", -- 0150
         x"c5",  x"cd",  x"4a",  x"02",  x"3e",  x"01",  x"cd",  x"03", -- 0158
         x"f0",  x"26",  x"cd",  x"51",  x"02",  x"af",  x"6c",  x"57", -- 0160
         x"67",  x"c1",  x"c3",  x"19",  x"c9",  x"83",  x"4c",  x"4f", -- 0168
         x"c3",  x"4d",  x"c1",  x"d8",  x"cd",  x"2c",  x"c9",  x"a0", -- 0170
         x"b7",  x"f9",  x"c0",  x"2c",  x"c9",  x"a1",  x"b7",  x"f9", -- 0178
         x"c0",  x"18",  x"cc",  x"86",  x"57",  x"49",  x"4e",  x"44", -- 0180
         x"4f",  x"d7",  x"6d",  x"c1",  x"d8",  x"cd",  x"56",  x"ce", -- 0188
         x"2c",  x"c9",  x"a0",  x"b7",  x"0b",  x"c1",  x"fa",  x"cc", -- 0190
         x"fa",  x"cc",  x"98",  x"cc",  x"2c",  x"c9",  x"20",  x"00", -- 0198
         x"7c",  x"d0",  x"2c",  x"c9",  x"05",  x"00",  x"51",  x"d1", -- 01A0
         x"2c",  x"c9",  x"9f",  x"b7",  x"f9",  x"c0",  x"2c",  x"c9", -- 01A8
         x"9d",  x"b7",  x"f9",  x"c0",  x"fa",  x"cc",  x"fa",  x"cc", -- 01B0
         x"98",  x"cc",  x"2c",  x"c9",  x"28",  x"00",  x"7c",  x"d0", -- 01B8
         x"2c",  x"c9",  x"05",  x"00",  x"51",  x"d1",  x"2c",  x"c9", -- 01C0
         x"9e",  x"b7",  x"f9",  x"c0",  x"2c",  x"c9",  x"9c",  x"b7", -- 01C8
         x"f9",  x"c0",  x"18",  x"cc",  x"83",  x"50",  x"49",  x"d8", -- 01D0
         x"83",  x"c1",  x"dc",  x"c1",  x"d1",  x"e1",  x"7c",  x"b7", -- 01D8
         x"28",  x"06",  x"7d",  x"e6",  x"c0",  x"b4",  x"e6",  x"fe", -- 01E0
         x"b2",  x"20",  x"1a",  x"cd",  x"4a",  x"02",  x"7b",  x"32", -- 01E8
         x"d5",  x"b7",  x"22",  x"d3",  x"b7",  x"cd",  x"51",  x"02", -- 01F0
         x"1e",  x"2f",  x"e1",  x"7d",  x"b4",  x"28",  x"01",  x"1c", -- 01F8
         x"cd",  x"0c",  x"f0",  x"18",  x"01",  x"e1",  x"c3",  x"1b", -- 0200
         x"c9",  x"83",  x"49",  x"4e",  x"cb",  x"d4",  x"c1",  x"11", -- 0208
         x"c2",  x"21",  x"a3",  x"b7",  x"d1",  x"cd",  x"4a",  x"02", -- 0210
         x"7b",  x"87",  x"87",  x"87",  x"e6",  x"7f",  x"57",  x"7e", -- 0218
         x"e6",  x"87",  x"b2",  x"77",  x"cd",  x"51",  x"02",  x"c3", -- 0220
         x"1b",  x"c9",  x"84",  x"49",  x"4e",  x"4b",  x"d0",  x"09", -- 0228
         x"c2",  x"33",  x"c2",  x"21",  x"d6",  x"b7",  x"18",  x"dc", -- 0230
         x"85",  x"42",  x"4c",  x"49",  x"4e",  x"cb",  x"2a",  x"c2", -- 0238
         x"42",  x"c2",  x"21",  x"a3",  x"b7",  x"cd",  x"4a",  x"02", -- 0240
         x"3e",  x"80",  x"ae",  x"77",  x"cd",  x"51",  x"02",  x"c3", -- 0248
         x"1b",  x"c9",  x"86",  x"42",  x"4c",  x"49",  x"4e",  x"4b", -- 0250
         x"d0",  x"38",  x"c2",  x"5d",  x"c2",  x"21",  x"d6",  x"b7", -- 0258
         x"18",  x"e3",  x"85",  x"50",  x"41",  x"50",  x"45",  x"d2", -- 0260
         x"52",  x"c2",  x"6c",  x"c2",  x"21",  x"a3",  x"b7",  x"cd", -- 0268
         x"4a",  x"02",  x"d1",  x"7b",  x"e6",  x"07",  x"57",  x"7e", -- 0270
         x"e6",  x"f8",  x"b2",  x"77",  x"cd",  x"51",  x"02",  x"c3", -- 0278
         x"1b",  x"c9",  x"85",  x"43",  x"4f",  x"4c",  x"4f",  x"d2", -- 0280
         x"62",  x"c2",  x"d8",  x"cd",  x"6a",  x"c2",  x"0f",  x"c2", -- 0288
         x"18",  x"cc",  x"85",  x"53",  x"4f",  x"55",  x"4e",  x"c4", -- 0290
         x"82",  x"c2",  x"9c",  x"c2",  x"d9",  x"21",  x"87",  x"b7", -- 0298
         x"06",  x"06",  x"cd",  x"4a",  x"02",  x"d1",  x"73",  x"2b", -- 02A0
         x"10",  x"fb",  x"1e",  x"35",  x"cd",  x"0c",  x"f0",  x"d9", -- 02A8
         x"c3",  x"1b",  x"c9",  x"83",  x"52",  x"2f",  x"d7",  x"92", -- 02B0
         x"c2",  x"bb",  x"c2",  x"e1",  x"7d",  x"fe",  x"05",  x"38", -- 02B8
         x"11",  x"db",  x"88",  x"e6",  x"9f",  x"d3",  x"88",  x"dd", -- 02C0
         x"e5",  x"e1",  x"7c",  x"1e",  x"31",  x"cd",  x"0c",  x"f0", -- 02C8
         x"18",  x"6c",  x"cd",  x"4a",  x"02",  x"7d",  x"d9",  x"fe", -- 02D0
         x"03",  x"30",  x"04",  x"1e",  x"02",  x"18",  x"02",  x"1e", -- 02D8
         x"0a",  x"16",  x"00",  x"2a",  x"b0",  x"b7",  x"19",  x"5e", -- 02E0
         x"23",  x"56",  x"eb",  x"f5",  x"cd",  x"51",  x"02",  x"f1", -- 02E8
         x"d1",  x"dd",  x"73",  x"05",  x"dd",  x"72",  x"06",  x"fe", -- 02F0
         x"03",  x"30",  x"25",  x"b7",  x"20",  x"09",  x"dd",  x"36", -- 02F8
         x"02",  x"00",  x"01",  x"00",  x"20",  x"18",  x"0b",  x"fe", -- 0300
         x"02",  x"20",  x"04",  x"dd",  x"36",  x"02",  x"fe",  x"01", -- 0308
         x"e0",  x"00",  x"db",  x"88",  x"f6",  x"60",  x"d3",  x"88", -- 0310
         x"11",  x"1d",  x"c3",  x"d5",  x"e9",  x"d9",  x"18",  x"1e", -- 0318
         x"fe",  x"03",  x"20",  x"08",  x"db",  x"88",  x"f6",  x"40", -- 0320
         x"e6",  x"df",  x"d3",  x"88",  x"11",  x"31",  x"c3",  x"d5", -- 0328
         x"e9",  x"d9",  x"16",  x"00",  x"dd",  x"5e",  x"02",  x"21", -- 0330
         x"00",  x"00",  x"ed",  x"6a",  x"d5",  x"e5",  x"c3",  x"1b", -- 0338
         x"c9",  x"85",  x"43",  x"4c",  x"4f",  x"41",  x"c4",  x"b3", -- 0340
         x"c2",  x"d8",  x"cd",  x"2c",  x"c9",  x"a4",  x"b7",  x"e0", -- 0348
         x"c0",  x"8a",  x"d0",  x"8a",  x"d0",  x"2c",  x"c9",  x"11", -- 0350
         x"00",  x"a5",  x"ca",  x"1b",  x"d5",  x"6e",  x"ce",  x"b9", -- 0358
         x"c2",  x"09",  x"cd",  x"5e",  x"ce",  x"2f",  x"d0",  x"e5", -- 0360
         x"ca",  x"68",  x"c9",  x"0a",  x"00",  x"09",  x"cd",  x"09", -- 0368
         x"cd",  x"56",  x"ce",  x"56",  x"ce",  x"68",  x"c9",  x"0a", -- 0370
         x"00",  x"34",  x"d3",  x"01",  x"2a",  x"50",  x"c9",  x"dc", -- 0378
         x"ff",  x"23",  x"cd",  x"68",  x"c9",  x"f0",  x"00",  x"fa", -- 0380
         x"ca",  x"1b",  x"d5",  x"2c",  x"c9",  x"0b",  x"00",  x"d3", -- 0388
         x"d2",  x"fa",  x"ca",  x"38",  x"cf",  x"64",  x"cd",  x"f8", -- 0390
         x"da",  x"02",  x"da",  x"d6",  x"cf",  x"cd",  x"cf",  x"95", -- 0398
         x"cd",  x"16",  x"cd",  x"5e",  x"ce",  x"ac",  x"d9",  x"23", -- 03A0
         x"cd",  x"77",  x"db",  x"8a",  x"d0",  x"04",  x"db",  x"96", -- 03A8
         x"d9",  x"f8",  x"da",  x"02",  x"da",  x"8a",  x"d0",  x"5e", -- 03B0
         x"ce",  x"2f",  x"d0",  x"f8",  x"da",  x"02",  x"da",  x"cb", -- 03B8
         x"c9",  x"5e",  x"ce",  x"cd",  x"cf",  x"3f",  x"cd",  x"56", -- 03C0
         x"ce",  x"6e",  x"ce",  x"56",  x"ce",  x"cb",  x"c9",  x"09", -- 03C8
         x"cd",  x"23",  x"cd",  x"2c",  x"c9",  x"04",  x"00",  x"b9", -- 03D0
         x"c2",  x"16",  x"cd",  x"23",  x"cd",  x"6e",  x"ce",  x"3f", -- 03D8
         x"de",  x"e5",  x"ca",  x"68",  x"c9",  x"0c",  x"00",  x"09", -- 03E0
         x"cd",  x"09",  x"cd",  x"56",  x"ce",  x"2c",  x"c9",  x"ff", -- 03E8
         x"00",  x"23",  x"cd",  x"2c",  x"c9",  x"ff",  x"00",  x"3d", -- 03F0
         x"d0",  x"68",  x"c9",  x"08",  x"00",  x"23",  x"cd",  x"cd", -- 03F8
         x"cf",  x"95",  x"cd",  x"cd",  x"cf",  x"64",  x"cd",  x"3d", -- 0400
         x"d0",  x"74",  x"cc",  x"68",  x"c9",  x"0c",  x"00",  x"34", -- 0408
         x"d3",  x"01",  x"2a",  x"09",  x"cd",  x"50",  x"c9",  x"ba", -- 0410
         x"ff",  x"23",  x"cd",  x"68",  x"c9",  x"0a",  x"00",  x"34", -- 0418
         x"d3",  x"01",  x"3f",  x"50",  x"c9",  x"08",  x"00",  x"2f", -- 0420
         x"cc",  x"34",  x"d3",  x"01",  x"3e",  x"7d",  x"c9",  x"a0", -- 0428
         x"ff",  x"68",  x"c9",  x"10",  x"00",  x"fa",  x"ca",  x"2c", -- 0430
         x"c9",  x"08",  x"00",  x"c7",  x"da",  x"cd",  x"cf",  x"6a", -- 0438
         x"de",  x"fa",  x"ca",  x"2c",  x"c9",  x"80",  x"00",  x"98", -- 0440
         x"cc",  x"cd",  x"cf",  x"64",  x"cd",  x"f8",  x"da",  x"31", -- 0448
         x"da",  x"5e",  x"ce",  x"3d",  x"d0",  x"68",  x"c9",  x"04", -- 0450
         x"00",  x"e3",  x"cf",  x"cd",  x"cf",  x"64",  x"cd",  x"2c", -- 0458
         x"c9",  x"ff",  x"00",  x"3d",  x"d0",  x"68",  x"c9",  x"04", -- 0460
         x"00",  x"2f",  x"cc",  x"7d",  x"c9",  x"54",  x"ff",  x"09", -- 0468
         x"cd",  x"50",  x"c9",  x"06",  x"00",  x"09",  x"cd",  x"09", -- 0470
         x"cd",  x"2c",  x"c9",  x"a4",  x"b7",  x"0b",  x"c1",  x"2c", -- 0478
         x"c9",  x"05",  x"00",  x"b9",  x"c2",  x"cd",  x"cf",  x"64", -- 0480
         x"cd",  x"2c",  x"c9",  x"ff",  x"00",  x"2f",  x"d0",  x"68", -- 0488
         x"c9",  x"0a",  x"00",  x"fa",  x"ca",  x"2c",  x"c9",  x"06", -- 0490
         x"00",  x"c7",  x"da",  x"18",  x"cc",  x"86",  x"56",  x"45", -- 0498
         x"52",  x"49",  x"46",  x"d9",  x"41",  x"c3",  x"d8",  x"cd", -- 04A0
         x"2c",  x"c9",  x"11",  x"00",  x"56",  x"ce",  x"49",  x"c0", -- 04A8
         x"18",  x"cc",  x"85",  x"43",  x"53",  x"41",  x"56",  x"c5", -- 04B0
         x"9d",  x"c4",  x"d8",  x"cd",  x"77",  x"ce",  x"2e",  x"d5", -- 04B8
         x"2c",  x"c9",  x"29",  x"20",  x"2c",  x"c9",  x"28",  x"46", -- 04C0
         x"f2",  x"cf",  x"2c",  x"c9",  x"09",  x"00",  x"98",  x"cc", -- 04C8
         x"b1",  x"cd",  x"f2",  x"cf",  x"2c",  x"c9",  x"0c",  x"00", -- 04D0
         x"98",  x"cc",  x"2c",  x"c9",  x"74",  x"00",  x"e3",  x"d4", -- 04D8
         x"f2",  x"cf",  x"d6",  x"cf",  x"56",  x"ce",  x"b9",  x"c2", -- 04E0
         x"04",  x"db",  x"96",  x"d9",  x"23",  x"cd",  x"8a",  x"d0", -- 04E8
         x"5e",  x"ce",  x"ac",  x"d9",  x"31",  x"cd",  x"2f",  x"d0", -- 04F0
         x"68",  x"c9",  x"3e",  x"00",  x"cb",  x"c9",  x"e7",  x"c9", -- 04F8
         x"77",  x"db",  x"f8",  x"da",  x"56",  x"ce",  x"cb",  x"c9", -- 0500
         x"23",  x"cd",  x"5e",  x"ce",  x"b9",  x"c2",  x"2c",  x"c9", -- 0508
         x"80",  x"00",  x"98",  x"cc",  x"e5",  x"ca",  x"68",  x"c9", -- 0510
         x"08",  x"00",  x"09",  x"cd",  x"56",  x"ce",  x"2f",  x"cc", -- 0518
         x"7d",  x"c9",  x"e6",  x"ff",  x"74",  x"cc",  x"68",  x"c9", -- 0520
         x"08",  x"00",  x"09",  x"cd",  x"56",  x"ce",  x"2f",  x"cc", -- 0528
         x"7d",  x"c9",  x"cc",  x"ff",  x"50",  x"c9",  x"06",  x"00", -- 0530
         x"09",  x"cd",  x"09",  x"cd",  x"a9",  x"d0",  x"68",  x"c9", -- 0538
         x"2a",  x"00",  x"77",  x"db",  x"6e",  x"ce",  x"56",  x"ce", -- 0540
         x"cb",  x"c9",  x"23",  x"cd",  x"5e",  x"ce",  x"b9",  x"c2", -- 0548
         x"2c",  x"c9",  x"80",  x"00",  x"98",  x"cc",  x"e5",  x"ca", -- 0550
         x"68",  x"c9",  x"08",  x"00",  x"09",  x"cd",  x"f2",  x"cf", -- 0558
         x"2f",  x"cc",  x"7d",  x"c9",  x"e6",  x"ff",  x"50",  x"c9", -- 0560
         x"04",  x"00",  x"f2",  x"cf",  x"66",  x"ce",  x"b9",  x"c2", -- 0568
         x"2c",  x"c9",  x"05",  x"00",  x"b9",  x"c2",  x"18",  x"cc", -- 0570
         x"84",  x"50",  x"4c",  x"4f",  x"d4",  x"b2",  x"c4",  x"81", -- 0578
         x"c5",  x"cd",  x"4a",  x"02",  x"d9",  x"3e",  x"30",  x"d1", -- 0580
         x"c1",  x"d9",  x"d1",  x"e1",  x"d9",  x"e1",  x"fd",  x"2b", -- 0588
         x"fd",  x"74",  x"00",  x"fd",  x"2b",  x"fd",  x"75",  x"00", -- 0590
         x"cb",  x"7a",  x"20",  x"04",  x"f6",  x"0a",  x"18",  x"07", -- 0598
         x"a7",  x"21",  x"00",  x"00",  x"ed",  x"52",  x"eb",  x"cb", -- 05A0
         x"78",  x"20",  x"04",  x"f6",  x"05",  x"18",  x"08",  x"a7", -- 05A8
         x"21",  x"00",  x"00",  x"ed",  x"42",  x"44",  x"4d",  x"60", -- 05B0
         x"69",  x"a7",  x"ed",  x"52",  x"38",  x"05",  x"c5",  x"e6", -- 05B8
         x"df",  x"18",  x"0a",  x"62",  x"6b",  x"a7",  x"ed",  x"42", -- 05C0
         x"d5",  x"e6",  x"ef",  x"59",  x"50",  x"4d",  x"44",  x"cb", -- 05C8
         x"3c",  x"cb",  x"1d",  x"d9",  x"08",  x"7c",  x"b7",  x"28", -- 05D0
         x"06",  x"7d",  x"e6",  x"c0",  x"b4",  x"e6",  x"fe",  x"b2", -- 05D8
         x"20",  x"17",  x"7b",  x"32",  x"d5",  x"b7",  x"22",  x"d3", -- 05E0
         x"b7",  x"d5",  x"1e",  x"30",  x"fd",  x"7e",  x"00",  x"fd", -- 05E8
         x"b6",  x"01",  x"20",  x"01",  x"1d",  x"cd",  x"09",  x"f0", -- 05F0
         x"d1",  x"08",  x"d9",  x"e3",  x"2b",  x"cb",  x"7c",  x"20", -- 05F8
         x"37",  x"e3",  x"a7",  x"ed",  x"52",  x"38",  x"1b",  x"d9", -- 0600
         x"cb",  x"67",  x"28",  x"08",  x"cb",  x"47",  x"28",  x"03", -- 0608
         x"23",  x"18",  x"01",  x"2b",  x"cb",  x"6f",  x"28",  x"1d", -- 0610
         x"cb",  x"4f",  x"28",  x"03",  x"13",  x"18",  x"16",  x"1b", -- 0618
         x"18",  x"13",  x"19",  x"09",  x"d9",  x"cb",  x"57",  x"28", -- 0620
         x"03",  x"23",  x"18",  x"01",  x"2b",  x"cb",  x"5f",  x"28", -- 0628
         x"03",  x"13",  x"18",  x"01",  x"1b",  x"d9",  x"18",  x"9b", -- 0630
         x"fd",  x"66",  x"01",  x"fd",  x"6e",  x"00",  x"e3",  x"fd", -- 0638
         x"23",  x"fd",  x"23",  x"d9",  x"e5",  x"d5",  x"cd",  x"51", -- 0640
         x"02",  x"c3",  x"1b",  x"c9",  x"84",  x"54",  x"45",  x"58", -- 0648
         x"d4",  x"74",  x"02",  x"d8",  x"cd",  x"f2",  x"cf",  x"81", -- 0650
         x"ce",  x"d6",  x"cf",  x"f4",  x"d4",  x"2e",  x"d5",  x"f2", -- 0658
         x"cf",  x"1b",  x"d5",  x"81",  x"ce",  x"d6",  x"cf",  x"13", -- 0660
         x"cb",  x"18",  x"cc",  x"84",  x"4c",  x"49",  x"4e",  x"c5", -- 0668
         x"4c",  x"c6",  x"d8",  x"cd",  x"23",  x"cd",  x"2c",  x"c9", -- 0670
         x"f0",  x"ff",  x"96",  x"cb",  x"2c",  x"c9",  x"17",  x"00", -- 0678
         x"51",  x"d1",  x"5f",  x"cf",  x"64",  x"cd",  x"83",  x"da", -- 0680
         x"09",  x"cd",  x"18",  x"cc",  x"85",  x"2d",  x"4d",  x"4f", -- 0688
         x"56",  x"c5",  x"6b",  x"c6",  x"d8",  x"cd",  x"72",  x"c6", -- 0690
         x"81",  x"ce",  x"13",  x"cb",  x"18",  x"cc",  x"81",  x"d2", -- 0698
         x"8c",  x"c6",  x"d8",  x"cd",  x"1b",  x"d5",  x"d6",  x"cf", -- 06A0
         x"16",  x"cd",  x"94",  x"c6",  x"18",  x"cc",  x"81",  x"d0", -- 06A8
         x"9e",  x"c6",  x"d8",  x"cd",  x"5e",  x"ce",  x"53",  x"c6", -- 06B0
         x"a2",  x"c6",  x"18",  x"cc",  x"81",  x"c8",  x"ae",  x"c6", -- 06B8
         x"d8",  x"cd",  x"72",  x"c6",  x"1b",  x"d5",  x"d6",  x"cf", -- 06C0
         x"81",  x"ce",  x"13",  x"cb",  x"18",  x"cc",  x"81",  x"d4", -- 06C8
         x"bc",  x"c6",  x"d8",  x"cd",  x"5f",  x"cf",  x"64",  x"cd", -- 06D0
         x"b3",  x"da",  x"18",  x"cc",  x"81",  x"c5",  x"ce",  x"c6", -- 06D8
         x"d8",  x"cd",  x"72",  x"c6",  x"81",  x"ce",  x"f4",  x"d4", -- 06E0
         x"18",  x"cc",  x"81",  x"cc",  x"dc",  x"c6",  x"d8",  x"cd", -- 06E8
         x"2c",  x"c9",  x"0c",  x"00",  x"a5",  x"ca",  x"5f",  x"cf", -- 06F0
         x"64",  x"cd",  x"e0",  x"de",  x"18",  x"cc",  x"81",  x"d3", -- 06F8
         x"ea",  x"c6",  x"d8",  x"cd",  x"2c",  x"c9",  x"0e",  x"00", -- 0700
         x"2c",  x"c9",  x"0f",  x"00",  x"8a",  x"d0",  x"cb",  x"c9", -- 0708
         x"23",  x"cd",  x"72",  x"c6",  x"fa",  x"cc",  x"d6",  x"cf", -- 0710
         x"94",  x"c6",  x"5e",  x"ce",  x"2f",  x"d0",  x"7d",  x"c9", -- 0718
         x"f0",  x"ff",  x"d6",  x"cf",  x"e0",  x"c6",  x"18",  x"cc", -- 0720
         x"81",  x"c4",  x"fe",  x"c6",  x"d8",  x"cd",  x"23",  x"cd", -- 0728
         x"c0",  x"c6",  x"2c",  x"c9",  x"10",  x"00",  x"16",  x"cd", -- 0730
         x"d6",  x"cf",  x"cb",  x"c9",  x"e7",  x"c9",  x"72",  x"c6", -- 0738
         x"e7",  x"c9",  x"5e",  x"ce",  x"2f",  x"d0",  x"94",  x"c6", -- 0740
         x"7d",  x"c9",  x"f2",  x"ff",  x"2c",  x"c9",  x"0f",  x"00", -- 0748
         x"e0",  x"c6",  x"18",  x"cc",  x"85",  x"43",  x"4c",  x"45", -- 0750
         x"41",  x"d2",  x"28",  x"c7",  x"d8",  x"cd",  x"5f",  x"cf", -- 0758
         x"95",  x"cd",  x"2c",  x"c9",  x"10",  x"00",  x"56",  x"ce", -- 0760
         x"cb",  x"c9",  x"e7",  x"c9",  x"e0",  x"c6",  x"7d",  x"c9", -- 0768
         x"fa",  x"ff",  x"18",  x"cc",  x"84",  x"4d",  x"4f",  x"56", -- 0770
         x"c5",  x"54",  x"c7",  x"d8",  x"cd",  x"2c",  x"c9",  x"10", -- 0778
         x"00",  x"56",  x"ce",  x"cb",  x"c9",  x"fa",  x"cc",  x"5f", -- 0780
         x"cf",  x"95",  x"cd",  x"e7",  x"c9",  x"72",  x"c6",  x"fa", -- 0788
         x"cc",  x"5f",  x"cf",  x"95",  x"cd",  x"e7",  x"c9",  x"94", -- 0790
         x"c6",  x"7d",  x"c9",  x"ea",  x"ff",  x"09",  x"cd",  x"09", -- 0798
         x"cd",  x"18",  x"cc",  x"84",  x"45",  x"44",  x"49",  x"d4", -- 07A0
         x"74",  x"c7",  x"d8",  x"cd",  x"5f",  x"cf",  x"95",  x"cd", -- 07A8
         x"2c",  x"c9",  x"a3",  x"b7",  x"cd",  x"c0",  x"2c",  x"c9", -- 07B0
         x"00",  x"00",  x"2c",  x"c9",  x"06",  x"00",  x"8a",  x"c2", -- 07B8
         x"56",  x"ce",  x"2c",  x"c9",  x"28",  x"00",  x"56",  x"ce", -- 07C0
         x"2c",  x"c9",  x"20",  x"00",  x"8c",  x"c1",  x"ee",  x"c6", -- 07C8
         x"2c",  x"c9",  x"07",  x"00",  x"6a",  x"c2",  x"2c",  x"c9", -- 07D0
         x"11",  x"00",  x"a5",  x"ca",  x"2c",  x"c9",  x"04",  x"00", -- 07D8
         x"2c",  x"c9",  x"20",  x"00",  x"66",  x"ce",  x"2c",  x"c9", -- 07E0
         x"10",  x"00",  x"8c",  x"c1",  x"c9",  x"ca",  x"23",  x"cd", -- 07E8
         x"23",  x"cd",  x"2c",  x"c9",  x"0c",  x"00",  x"3d",  x"d0", -- 07F0
         x"68",  x"c9",  x"20",  x"00",  x"a5",  x"ca",  x"2c",  x"c9", -- 07F8
         x"10",  x"00",  x"56",  x"ce",  x"cb",  x"c9",  x"e7",  x"c9", -- 0800
         x"56",  x"ce",  x"73",  x"c1",  x"e7",  x"c9",  x"d2",  x"c6", -- 0808
         x"7d",  x"c9",  x"f4",  x"ff",  x"fa",  x"ca",  x"50",  x"c9", -- 0810
         x"16",  x"00",  x"23",  x"cd",  x"2c",  x"c9",  x"0d",  x"00", -- 0818
         x"3d",  x"d0",  x"68",  x"c9",  x"08",  x"00",  x"2c",  x"c9", -- 0820
         x"0a",  x"00",  x"a5",  x"ca",  x"a5",  x"ca",  x"2c",  x"c9", -- 0828
         x"13",  x"00",  x"3d",  x"d0",  x"68",  x"c9",  x"b6",  x"ff", -- 0830
         x"2c",  x"c9",  x"10",  x"00",  x"56",  x"ce",  x"cb",  x"c9", -- 0838
         x"2c",  x"c9",  x"54",  x"b2",  x"e7",  x"c9",  x"2c",  x"c9", -- 0840
         x"28",  x"00",  x"02",  x"da",  x"98",  x"cc",  x"e7",  x"c9", -- 0848
         x"72",  x"c6",  x"81",  x"ce",  x"56",  x"ce",  x"cb",  x"c9", -- 0850
         x"45",  x"cc",  x"23",  x"cd",  x"cd",  x"c0",  x"a9",  x"d0", -- 0858
         x"68",  x"c9",  x"06",  x"00",  x"50",  x"c9",  x"04",  x"00", -- 0860
         x"77",  x"ce",  x"6d",  x"cc",  x"a4",  x"cd",  x"d6",  x"cf", -- 0868
         x"5a",  x"cc",  x"d6",  x"cf",  x"7d",  x"c9",  x"e2",  x"ff", -- 0870
         x"09",  x"cd",  x"09",  x"cd",  x"7d",  x"c9",  x"c2",  x"ff", -- 0878
         x"56",  x"ce",  x"2c",  x"c9",  x"28",  x"00",  x"56",  x"ce", -- 0880
         x"2c",  x"c9",  x"20",  x"00",  x"8c",  x"c1",  x"2c",  x"c9", -- 0888
         x"12",  x"00",  x"a5",  x"ca",  x"2c",  x"c9",  x"12",  x"00", -- 0890
         x"56",  x"ce",  x"73",  x"c1",  x"2c",  x"c9",  x"a3",  x"b7", -- 0898
         x"f9",  x"c0",  x"18",  x"cc",  x"84",  x"44",  x"55",  x"4d", -- 08A0
         x"d0",  x"78",  x"c5",  x"ad",  x"c8",  x"1e",  x"2c",  x"cd", -- 08A8
         x"0c",  x"f0",  x"cd",  x"0c",  x"f0",  x"d1",  x"e1",  x"c5", -- 08B0
         x"42",  x"4b",  x"0b",  x"78",  x"07",  x"38",  x"4d",  x"1e", -- 08B8
         x"1a",  x"cd",  x"0c",  x"f0",  x"16",  x"08",  x"1e",  x"2b", -- 08C0
         x"cd",  x"0c",  x"f0",  x"7e",  x"1e",  x"1c",  x"cd",  x"0c", -- 08C8
         x"f0",  x"23",  x"15",  x"20",  x"f1",  x"11",  x"f8",  x"ff", -- 08D0
         x"19",  x"3e",  x"09",  x"1e",  x"24",  x"cd",  x"0c",  x"f0", -- 08D8
         x"16",  x"08",  x"7e",  x"e6",  x"7f",  x"fe",  x"20",  x"30", -- 08E0
         x"02",  x"3e",  x"2e",  x"1e",  x"24",  x"cd",  x"0c",  x"f0", -- 08E8
         x"23",  x"0b",  x"15",  x"20",  x"ed",  x"1e",  x"24",  x"3e", -- 08F0
         x"0d",  x"cd",  x"0c",  x"f0",  x"3e",  x"0a",  x"cd",  x"0c", -- 08F8
         x"f0",  x"1e",  x"0e",  x"cd",  x"0c",  x"f0",  x"30",  x"02", -- 0900
         x"06",  x"ff",  x"18",  x"af",  x"c1",  x"c3",  x"1b",  x"c9", -- 0908
         x"84",  x"54",  x"41",  x"53",  x"cb",  x"a4",  x"c8",  x"1b", -- 0910
         x"c9",  x"d5",  x"e5",  x"0a",  x"03",  x"6f",  x"0a",  x"03", -- 0918
         x"67",  x"5e",  x"23",  x"56",  x"eb",  x"e9",  x"83",  x"4c", -- 0920
         x"49",  x"d4",  x"00",  x"00",  x"2e",  x"c9",  x"0a",  x"03", -- 0928
         x"6f",  x"0a",  x"03",  x"67",  x"c3",  x"1a",  x"c9",  x"87", -- 0930
         x"45",  x"58",  x"45",  x"43",  x"55",  x"54",  x"c5",  x"26", -- 0938
         x"c9",  x"43",  x"c9",  x"e1",  x"c3",  x"21",  x"c9",  x"86", -- 0940
         x"42",  x"52",  x"41",  x"4e",  x"43",  x"c8",  x"37",  x"c9", -- 0948
         x"52",  x"c9",  x"60",  x"69",  x"5e",  x"23",  x"56",  x"2b", -- 0950
         x"19",  x"4d",  x"44",  x"c3",  x"1b",  x"c9",  x"87",  x"30", -- 0958
         x"42",  x"52",  x"41",  x"4e",  x"43",  x"c8",  x"47",  x"c9", -- 0960
         x"6a",  x"c9",  x"e1",  x"7d",  x"b4",  x"28",  x"e3",  x"03", -- 0968
         x"03",  x"c3",  x"1b",  x"c9",  x"86",  x"28",  x"4c",  x"4f", -- 0970
         x"4f",  x"50",  x"a9",  x"5e",  x"c9",  x"7f",  x"c9",  x"11", -- 0978
         x"01",  x"00",  x"fd",  x"7e",  x"00",  x"83",  x"fd",  x"77", -- 0980
         x"00",  x"5f",  x"fd",  x"7e",  x"01",  x"8a",  x"fd",  x"77", -- 0988
         x"01",  x"cb",  x"12",  x"57",  x"38",  x"0a",  x"7b",  x"fd", -- 0990
         x"96",  x"02",  x"7a",  x"fd",  x"9e",  x"03",  x"18",  x"08", -- 0998
         x"fd",  x"7e",  x"02",  x"93",  x"fd",  x"7e",  x"03",  x"9a", -- 09A0
         x"07",  x"38",  x"a7",  x"11",  x"04",  x"00",  x"fd",  x"19", -- 09A8
         x"03",  x"03",  x"c3",  x"1b",  x"c9",  x"87",  x"28",  x"2b", -- 09B0
         x"4c",  x"4f",  x"4f",  x"50",  x"a9",  x"74",  x"c9",  x"c1", -- 09B8
         x"c9",  x"d1",  x"18",  x"be",  x"84",  x"28",  x"44",  x"4f", -- 09C0
         x"a9",  x"b5",  x"c9",  x"cd",  x"c9",  x"11",  x"fc",  x"ff", -- 09C8
         x"fd",  x"19",  x"d1",  x"fd",  x"73",  x"00",  x"fd",  x"72", -- 09D0
         x"01",  x"d1",  x"fd",  x"73",  x"02",  x"fd",  x"72",  x"03", -- 09D8
         x"c3",  x"1b",  x"c9",  x"81",  x"c9",  x"c4",  x"c9",  x"e9", -- 09E0
         x"c9",  x"fd",  x"6e",  x"00",  x"fd",  x"66",  x"01",  x"c3", -- 09E8
         x"1a",  x"c9",  x"85",  x"44",  x"49",  x"47",  x"49",  x"d4", -- 09F0
         x"e3",  x"c9",  x"fc",  x"c9",  x"e1",  x"d1",  x"7b",  x"d6", -- 09F8
         x"30",  x"38",  x"13",  x"fe",  x"0a",  x"38",  x"06",  x"d6", -- 0A00
         x"07",  x"fe",  x"0a",  x"38",  x"09",  x"bd",  x"30",  x"06", -- 0A08
         x"5f",  x"2e",  x"01",  x"d5",  x"18",  x"01",  x"6c",  x"c3", -- 0A10
         x"1a",  x"c9",  x"86",  x"28",  x"46",  x"49",  x"4e",  x"44", -- 0A18
         x"a9",  x"f2",  x"c9",  x"25",  x"ca",  x"d1",  x"e1",  x"e5", -- 0A20
         x"1a",  x"ae",  x"e6",  x"3f",  x"20",  x"1f",  x"23",  x"13", -- 0A28
         x"1a",  x"ae",  x"87",  x"20",  x"16",  x"30",  x"f7",  x"21", -- 0A30
         x"05",  x"00",  x"19",  x"e3",  x"1b",  x"1a",  x"cb",  x"7f", -- 0A38
         x"28",  x"fa",  x"5f",  x"16",  x"00",  x"21",  x"01",  x"00", -- 0A40
         x"d5",  x"18",  x"15",  x"38",  x"06",  x"13",  x"1a",  x"cb", -- 0A48
         x"7f",  x"28",  x"fa",  x"13",  x"eb",  x"5e",  x"23",  x"56", -- 0A50
         x"7b",  x"b2",  x"20",  x"ca",  x"e1",  x"21",  x"00",  x"00", -- 0A58
         x"c3",  x"1a",  x"c9",  x"87",  x"45",  x"4e",  x"43",  x"4c", -- 0A60
         x"4f",  x"53",  x"c5",  x"1a",  x"ca",  x"6f",  x"ca",  x"d1", -- 0A68
         x"e1",  x"e5",  x"08",  x"7b",  x"11",  x"ff",  x"ff",  x"2b", -- 0A70
         x"23",  x"13",  x"be",  x"28",  x"fb",  x"d5",  x"08",  x"7e", -- 0A78
         x"b7",  x"20",  x"06",  x"13",  x"d5",  x"1b",  x"d5",  x"18", -- 0A80
         x"12",  x"08",  x"23",  x"13",  x"be",  x"28",  x"09",  x"08", -- 0A88
         x"7e",  x"b7",  x"20",  x"f5",  x"d5",  x"d5",  x"18",  x"03", -- 0A90
         x"d5",  x"13",  x"d5",  x"c3",  x"1b",  x"c9",  x"84",  x"45", -- 0A98
         x"4d",  x"49",  x"d4",  x"63",  x"ca",  x"d8",  x"cd",  x"b5", -- 0AA0
         x"ca",  x"5e",  x"ce",  x"55",  x"cf",  x"3f",  x"cd",  x"18", -- 0AA8
         x"cc",  x"81",  x"a0",  x"9e",  x"ca",  x"b7",  x"ca",  x"e1", -- 0AB0
         x"7d",  x"e6",  x"7f",  x"1e",  x"24",  x"cd",  x"0c",  x"f0", -- 0AB8
         x"c3",  x"1b",  x"c9",  x"83",  x"4b",  x"45",  x"d9",  x"b1", -- 0AC0
         x"ca",  x"cb",  x"ca",  x"1e",  x"16",  x"cd",  x"0c",  x"f0", -- 0AC8
         x"b7",  x"28",  x"f8",  x"6f",  x"26",  x"00",  x"c3",  x"1a", -- 0AD0
         x"c9",  x"89",  x"3f",  x"54",  x"45",  x"52",  x"4d",  x"49", -- 0AD8
         x"4e",  x"41",  x"cc",  x"c3",  x"ca",  x"e7",  x"ca",  x"21", -- 0AE0
         x"00",  x"00",  x"1e",  x"0e",  x"cd",  x"0c",  x"f0",  x"30", -- 0AE8
         x"01",  x"23",  x"c3",  x"1a",  x"c9",  x"82",  x"43",  x"d2", -- 0AF0
         x"d9",  x"ca",  x"fc",  x"ca",  x"1e",  x"24",  x"3e",  x"0a", -- 0AF8
         x"cd",  x"0c",  x"f0",  x"3e",  x"0d",  x"cd",  x"0c",  x"f0", -- 0B00
         x"c3",  x"1b",  x"c9",  x"85",  x"43",  x"4d",  x"4f",  x"56", -- 0B08
         x"c5",  x"f5",  x"ca",  x"15",  x"cb",  x"d9",  x"c1",  x"d1", -- 0B10
         x"e1",  x"78",  x"b1",  x"28",  x"02",  x"ed",  x"b0",  x"d9", -- 0B18
         x"c3",  x"1b",  x"c9",  x"82",  x"55",  x"aa",  x"0b",  x"cb", -- 0B20
         x"2a",  x"cb",  x"e1",  x"d9",  x"c1",  x"11",  x"00",  x"00", -- 0B28
         x"63",  x"6b",  x"d9",  x"16",  x"10",  x"d9",  x"29",  x"cb", -- 0B30
         x"13",  x"cb",  x"12",  x"d9",  x"29",  x"30",  x"06",  x"d9", -- 0B38
         x"09",  x"30",  x"01",  x"13",  x"d9",  x"15",  x"20",  x"ed", -- 0B40
         x"d9",  x"e5",  x"d5",  x"d9",  x"c3",  x"1b",  x"c9",  x"82", -- 0B48
         x"55",  x"af",  x"23",  x"cb",  x"56",  x"cb",  x"21",  x"05", -- 0B50
         x"00",  x"39",  x"56",  x"70",  x"2b",  x"5e",  x"71",  x"c1", -- 0B58
         x"e1",  x"7d",  x"91",  x"7c",  x"98",  x"38",  x"07",  x"21", -- 0B60
         x"ff",  x"ff",  x"54",  x"5c",  x"18",  x"1c",  x"3e",  x"10", -- 0B68
         x"a7",  x"cb",  x"13",  x"cb",  x"12",  x"cb",  x"15",  x"cb", -- 0B70
         x"14",  x"30",  x"05",  x"a7",  x"ed",  x"42",  x"18",  x"06", -- 0B78
         x"ed",  x"42",  x"30",  x"02",  x"09",  x"1b",  x"13",  x"3d", -- 0B80
         x"20",  x"e6",  x"c1",  x"e5",  x"d5",  x"c3",  x"1b",  x"c9", -- 0B88
         x"83",  x"41",  x"4e",  x"c4",  x"4f",  x"cb",  x"98",  x"cb", -- 0B90
         x"e1",  x"d1",  x"7d",  x"a3",  x"6f",  x"7c",  x"a2",  x"67", -- 0B98
         x"c3",  x"1a",  x"c9",  x"82",  x"4f",  x"d2",  x"90",  x"cb", -- 0BA0
         x"aa",  x"cb",  x"e1",  x"d1",  x"7d",  x"b3",  x"6f",  x"7c", -- 0BA8
         x"b2",  x"67",  x"c3",  x"1a",  x"c9",  x"83",  x"58",  x"4f", -- 0BB0
         x"d2",  x"a3",  x"cb",  x"bd",  x"cb",  x"e1",  x"d1",  x"7d", -- 0BB8
         x"ab",  x"6f",  x"7c",  x"aa",  x"67",  x"c3",  x"1a",  x"c9", -- 0BC0
         x"83",  x"53",  x"50",  x"c0",  x"b5",  x"cb",  x"d0",  x"cb", -- 0BC8
         x"21",  x"00",  x"00",  x"39",  x"c3",  x"1a",  x"c9",  x"83", -- 0BD0
         x"53",  x"50",  x"a1",  x"c8",  x"cb",  x"df",  x"cb",  x"2a", -- 0BD8
         x"7e",  x"01",  x"11",  x"06",  x"00",  x"19",  x"5e",  x"23", -- 0BE0
         x"56",  x"eb",  x"f9",  x"c3",  x"1b",  x"c9",  x"83",  x"52", -- 0BE8
         x"50",  x"c0",  x"d7",  x"cb",  x"f6",  x"cb",  x"fd",  x"e5", -- 0BF0
         x"c3",  x"1b",  x"c9",  x"83",  x"52",  x"50",  x"a1",  x"ee", -- 0BF8
         x"cb",  x"03",  x"cc",  x"2a",  x"7e",  x"01",  x"11",  x"08", -- 0C00
         x"00",  x"19",  x"5e",  x"23",  x"56",  x"d5",  x"fd",  x"e1", -- 0C08
         x"c3",  x"1b",  x"c9",  x"82",  x"3b",  x"d3",  x"fb",  x"cb", -- 0C10
         x"1a",  x"cc",  x"fd",  x"4e",  x"00",  x"fd",  x"23",  x"fd", -- 0C18
         x"46",  x"00",  x"fd",  x"23",  x"c3",  x"1b",  x"c9",  x"85", -- 0C20
         x"4c",  x"45",  x"41",  x"56",  x"c5",  x"13",  x"cc",  x"31", -- 0C28
         x"cc",  x"fd",  x"7e",  x"00",  x"fd",  x"77",  x"02",  x"fd", -- 0C30
         x"7e",  x"01",  x"fd",  x"77",  x"03",  x"c3",  x"1b",  x"c9", -- 0C38
         x"82",  x"3e",  x"d2",  x"27",  x"cc",  x"47",  x"cc",  x"fd", -- 0C40
         x"2b",  x"fd",  x"2b",  x"d1",  x"fd",  x"73",  x"00",  x"fd", -- 0C48
         x"72",  x"01",  x"c3",  x"1b",  x"c9",  x"82",  x"52",  x"be", -- 0C50
         x"40",  x"cc",  x"5c",  x"cc",  x"fd",  x"6e",  x"00",  x"fd", -- 0C58
         x"23",  x"fd",  x"66",  x"00",  x"fd",  x"23",  x"c3",  x"1a", -- 0C60
         x"c9",  x"81",  x"d2",  x"55",  x"cc",  x"e9",  x"c9",  x"82", -- 0C68
         x"30",  x"bd",  x"69",  x"cc",  x"76",  x"cc",  x"e1",  x"7c", -- 0C70
         x"b5",  x"21",  x"00",  x"00",  x"20",  x"01",  x"23",  x"c3", -- 0C78
         x"1a",  x"c9",  x"82",  x"30",  x"bc",  x"6f",  x"cc",  x"89", -- 0C80
         x"cc",  x"e1",  x"29",  x"21",  x"00",  x"00",  x"30",  x"01", -- 0C88
         x"23",  x"c3",  x"1a",  x"c9",  x"81",  x"ab",  x"82",  x"cc", -- 0C90
         x"9a",  x"cc",  x"d1",  x"e1",  x"19",  x"c3",  x"1a",  x"c9", -- 0C98
         x"82",  x"44",  x"ab",  x"94",  x"cc",  x"a7",  x"cc",  x"21", -- 0CA0
         x"06",  x"00",  x"39",  x"5e",  x"71",  x"23",  x"56",  x"70", -- 0CA8
         x"c1",  x"e1",  x"19",  x"eb",  x"e1",  x"7d",  x"89",  x"6f", -- 0CB0
         x"7c",  x"88",  x"67",  x"c1",  x"d5",  x"c3",  x"1a",  x"c9", -- 0CB8
         x"85",  x"4d",  x"49",  x"4e",  x"55",  x"d3",  x"a0",  x"cc", -- 0CC0
         x"ca",  x"cc",  x"21",  x"00",  x"00",  x"d1",  x"b7",  x"ed", -- 0CC8
         x"52",  x"c3",  x"1a",  x"c9",  x"86",  x"44",  x"4d",  x"49", -- 0CD0
         x"4e",  x"55",  x"d3",  x"c0",  x"cc",  x"df",  x"cc",  x"e1", -- 0CD8
         x"d1",  x"af",  x"93",  x"5f",  x"3e",  x"00",  x"9a",  x"57", -- 0CE0
         x"3e",  x"00",  x"9d",  x"6f",  x"3e",  x"00",  x"9c",  x"67", -- 0CE8
         x"c3",  x"19",  x"c9",  x"84",  x"4f",  x"56",  x"45",  x"d2", -- 0CF0
         x"d4",  x"cc",  x"fc",  x"cc",  x"d1",  x"e1",  x"e5",  x"c3", -- 0CF8
         x"19",  x"c9",  x"84",  x"44",  x"52",  x"4f",  x"d0",  x"f3", -- 0D00
         x"cc",  x"0b",  x"cd",  x"e1",  x"c3",  x"1b",  x"c9",  x"84", -- 0D08
         x"53",  x"57",  x"41",  x"d0",  x"02",  x"cd",  x"18",  x"cd", -- 0D10
         x"e1",  x"e3",  x"c3",  x"1a",  x"c9",  x"83",  x"44",  x"55", -- 0D18
         x"d0",  x"0f",  x"cd",  x"25",  x"cd",  x"e1",  x"e5",  x"c3", -- 0D20
         x"1a",  x"c9",  x"84",  x"32",  x"44",  x"55",  x"d0",  x"1d", -- 0D28
         x"cd",  x"33",  x"cd",  x"e1",  x"d1",  x"d5",  x"e5",  x"c3", -- 0D30
         x"19",  x"c9",  x"82",  x"2b",  x"a1",  x"2a",  x"cd",  x"41", -- 0D38
         x"cd",  x"e1",  x"d1",  x"7e",  x"83",  x"77",  x"23",  x"7e", -- 0D40
         x"8a",  x"77",  x"c3",  x"1b",  x"c9",  x"86",  x"54",  x"4f", -- 0D48
         x"47",  x"47",  x"4c",  x"c5",  x"3a",  x"cd",  x"58",  x"cd", -- 0D50
         x"d1",  x"e1",  x"7e",  x"ab",  x"77",  x"c3",  x"1b",  x"c9", -- 0D58
         x"81",  x"c0",  x"4d",  x"cd",  x"66",  x"cd",  x"e1",  x"5e", -- 0D60
         x"23",  x"56",  x"d5",  x"c3",  x"1b",  x"c9",  x"82",  x"43", -- 0D68
         x"c0",  x"60",  x"cd",  x"75",  x"cd",  x"e1",  x"6e",  x"26", -- 0D70
         x"00",  x"c3",  x"1a",  x"c9",  x"82",  x"32",  x"c0",  x"6e", -- 0D78
         x"cd",  x"83",  x"cd",  x"e1",  x"5e",  x"23",  x"56",  x"23", -- 0D80
         x"7e",  x"23",  x"66",  x"6f",  x"e5",  x"d5",  x"c3",  x"1b", -- 0D88
         x"c9",  x"81",  x"a1",  x"7c",  x"cd",  x"97",  x"cd",  x"e1", -- 0D90
         x"d1",  x"73",  x"23",  x"72",  x"c3",  x"1b",  x"c9",  x"82", -- 0D98
         x"43",  x"a1",  x"91",  x"cd",  x"a6",  x"cd",  x"e1",  x"d1", -- 0DA0
         x"73",  x"c3",  x"1b",  x"c9",  x"82",  x"32",  x"a1",  x"9f", -- 0DA8
         x"cd",  x"b3",  x"cd",  x"e1",  x"d1",  x"73",  x"23",  x"72", -- 0DB0
         x"23",  x"d1",  x"73",  x"23",  x"72",  x"c3",  x"1b",  x"c9", -- 0DB8
         x"c1",  x"ba",  x"ac",  x"cd",  x"d8",  x"cd",  x"83",  x"d1", -- 0DC0
         x"3e",  x"d1",  x"7b",  x"cf",  x"64",  x"cd",  x"6d",  x"cf", -- 0DC8
         x"95",  x"cd",  x"b8",  x"d6",  x"0a",  x"d2",  x"5d",  x"d2", -- 0DD0
         x"fd",  x"2b",  x"fd",  x"70",  x"00",  x"fd",  x"2b",  x"fd", -- 0DD8
         x"71",  x"00",  x"13",  x"4b",  x"42",  x"c3",  x"1b",  x"c9", -- 0DE0
         x"c1",  x"bb",  x"c0",  x"cd",  x"d8",  x"cd",  x"ad",  x"d1", -- 0DE8
         x"e4",  x"d1",  x"18",  x"cc",  x"1f",  x"d2",  x"fb",  x"d1", -- 0DF0
         x"18",  x"cc",  x"88",  x"43",  x"4f",  x"4e",  x"53",  x"54", -- 0DF8
         x"41",  x"4e",  x"d4",  x"e8",  x"cd",  x"d8",  x"cd",  x"b8", -- 0E00
         x"d6",  x"1f",  x"d2",  x"0e",  x"d0",  x"5d",  x"d2",  x"13", -- 0E08
         x"eb",  x"5e",  x"23",  x"56",  x"d5",  x"c3",  x"1b",  x"c9", -- 0E10
         x"88",  x"56",  x"41",  x"52",  x"49",  x"41",  x"42",  x"4c", -- 0E18
         x"c5",  x"fa",  x"cd",  x"d8",  x"cd",  x"05",  x"ce",  x"5d", -- 0E20
         x"d2",  x"13",  x"d5",  x"c3",  x"1b",  x"c9",  x"84",  x"55", -- 0E28
         x"53",  x"45",  x"d2",  x"18",  x"ce",  x"d8",  x"cd",  x"05", -- 0E30
         x"ce",  x"5d",  x"d2",  x"13",  x"eb",  x"5e",  x"23",  x"56", -- 0E38
         x"2a",  x"7e",  x"01",  x"19",  x"c3",  x"1a",  x"c9",  x"84", -- 0E40
         x"4e",  x"45",  x"58",  x"d4",  x"2e",  x"ce",  x"0f",  x"ce", -- 0E48
         x"1b",  x"c9",  x"81",  x"b0",  x"47",  x"ce",  x"0f",  x"ce", -- 0E50
         x"00",  x"00",  x"81",  x"b1",  x"52",  x"ce",  x"0f",  x"ce", -- 0E58
         x"01",  x"00",  x"81",  x"b2",  x"5a",  x"ce",  x"0f",  x"ce", -- 0E60
         x"02",  x"00",  x"81",  x"b3",  x"62",  x"ce",  x"0f",  x"ce", -- 0E68
         x"03",  x"00",  x"82",  x"42",  x"cc",  x"6a",  x"ce",  x"0f", -- 0E70
         x"ce",  x"20",  x"00",  x"83",  x"43",  x"2f",  x"cc",  x"72", -- 0E78
         x"ce",  x"0f",  x"ce",  x"20",  x"00",  x"85",  x"42",  x"2f", -- 0E80
         x"42",  x"55",  x"c6",  x"7b",  x"ce",  x"0f",  x"ce",  x"00", -- 0E88
         x"02",  x"85",  x"42",  x"2f",  x"53",  x"43",  x"d2",  x"85", -- 0E90
         x"ce",  x"0f",  x"ce",  x"01",  x"00",  x"87",  x"2b",  x"4f", -- 0E98
         x"52",  x"49",  x"47",  x"49",  x"ce",  x"91",  x"ce",  x"d8", -- 0EA0
         x"cd",  x"2c",  x"c9",  x"18",  x"c0",  x"98",  x"cc",  x"18", -- 0EA8
         x"cc",  x"82",  x"53",  x"b0",  x"9d",  x"ce",  x"3b",  x"ce", -- 0EB0
         x"06",  x"00",  x"82",  x"52",  x"b0",  x"b1",  x"ce",  x"3b", -- 0EB8
         x"ce",  x"08",  x"00",  x"83",  x"54",  x"49",  x"c2",  x"ba", -- 0EC0
         x"ce",  x"3b",  x"ce",  x"0a",  x"00",  x"85",  x"57",  x"49", -- 0EC8
         x"44",  x"54",  x"c8",  x"c3",  x"ce",  x"3b",  x"ce",  x"0c", -- 0ED0
         x"00",  x"87",  x"57",  x"41",  x"52",  x"4e",  x"49",  x"4e", -- 0ED8
         x"c7",  x"cd",  x"ce",  x"3b",  x"ce",  x"0e",  x"00",  x"85", -- 0EE0
         x"46",  x"45",  x"4e",  x"43",  x"c5",  x"d9",  x"ce",  x"3b", -- 0EE8
         x"ce",  x"10",  x"00",  x"82",  x"44",  x"d0",  x"e7",  x"ce", -- 0EF0
         x"3b",  x"ce",  x"12",  x"00",  x"88",  x"56",  x"4f",  x"43", -- 0EF8
         x"2d",  x"4c",  x"49",  x"4e",  x"cb",  x"f3",  x"ce",  x"3b", -- 0F00
         x"ce",  x"14",  x"00",  x"85",  x"46",  x"49",  x"52",  x"53", -- 0F08
         x"d4",  x"fc",  x"ce",  x"3b",  x"ce",  x"16",  x"00",  x"85", -- 0F10
         x"4c",  x"49",  x"4d",  x"49",  x"d4",  x"0b",  x"cf",  x"3b", -- 0F18
         x"ce",  x"18",  x"00",  x"85",  x"49",  x"4f",  x"54",  x"41", -- 0F20
         x"c2",  x"17",  x"cf",  x"3b",  x"ce",  x"1a",  x"00",  x"86", -- 0F28
         x"4f",  x"46",  x"46",  x"53",  x"45",  x"d4",  x"23",  x"cf", -- 0F30
         x"3b",  x"ce",  x"1c",  x"00",  x"83",  x"42",  x"4c",  x"cb", -- 0F38
         x"2f",  x"cf",  x"3b",  x"ce",  x"1e",  x"00",  x"82",  x"49", -- 0F40
         x"ce",  x"3c",  x"cf",  x"3b",  x"ce",  x"20",  x"00",  x"83", -- 0F48
         x"4f",  x"55",  x"d4",  x"46",  x"cf",  x"3b",  x"ce",  x"22", -- 0F50
         x"00",  x"83",  x"53",  x"43",  x"d2",  x"4f",  x"cf",  x"3b", -- 0F58
         x"ce",  x"24",  x"00",  x"87",  x"43",  x"4f",  x"4e",  x"54", -- 0F60
         x"45",  x"58",  x"d4",  x"59",  x"cf",  x"3b",  x"ce",  x"26", -- 0F68
         x"00",  x"87",  x"43",  x"55",  x"52",  x"52",  x"45",  x"4e", -- 0F70
         x"d4",  x"63",  x"cf",  x"3b",  x"ce",  x"28",  x"00",  x"85", -- 0F78
         x"53",  x"54",  x"41",  x"54",  x"c5",  x"71",  x"cf",  x"3b", -- 0F80
         x"ce",  x"2a",  x"00",  x"84",  x"42",  x"41",  x"53",  x"c5", -- 0F88
         x"7f",  x"cf",  x"3b",  x"ce",  x"2c",  x"00",  x"83",  x"44", -- 0F90
         x"50",  x"cc",  x"8b",  x"cf",  x"3b",  x"ce",  x"2e",  x"00", -- 0F98
         x"83",  x"46",  x"4c",  x"c4",  x"96",  x"cf",  x"3b",  x"ce", -- 0FA0
         x"30",  x"00",  x"83",  x"43",  x"53",  x"d0",  x"a0",  x"cf", -- 0FA8
         x"3b",  x"ce",  x"32",  x"00",  x"82",  x"52",  x"a3",  x"aa", -- 0FB0
         x"cf",  x"3b",  x"ce",  x"34",  x"00",  x"83",  x"48",  x"4c", -- 0FB8
         x"c4",  x"b4",  x"cf",  x"3b",  x"ce",  x"36",  x"00",  x"83", -- 0FC0
         x"52",  x"45",  x"c3",  x"bd",  x"cf",  x"3b",  x"ce",  x"38", -- 0FC8
         x"00",  x"82",  x"31",  x"ab",  x"c7",  x"cf",  x"d8",  x"cd", -- 0FD0
         x"5e",  x"ce",  x"98",  x"cc",  x"18",  x"cc",  x"82",  x"32", -- 0FD8
         x"ab",  x"d1",  x"cf",  x"d8",  x"cd",  x"66",  x"ce",  x"98", -- 0FE0
         x"cc",  x"18",  x"cc",  x"84",  x"48",  x"45",  x"52",  x"c5", -- 0FE8
         x"de",  x"cf",  x"d8",  x"cd",  x"f8",  x"ce",  x"64",  x"cd", -- 0FF0
         x"18",  x"cc",  x"85",  x"41",  x"4c",  x"4c",  x"4f",  x"d4", -- 0FF8
         x"eb",  x"cf",  x"d8",  x"cd",  x"f8",  x"ce",  x"3f",  x"cd", -- 1000
         x"18",  x"cc",  x"81",  x"ac",  x"fa",  x"cf",  x"d8",  x"cd", -- 1008
         x"f2",  x"cf",  x"66",  x"ce",  x"02",  x"d0",  x"95",  x"cd", -- 1010
         x"18",  x"cc",  x"82",  x"43",  x"ac",  x"0a",  x"d0",  x"d8", -- 1018
         x"cd",  x"f2",  x"cf",  x"5e",  x"ce",  x"02",  x"d0",  x"a4", -- 1020
         x"cd",  x"18",  x"cc",  x"81",  x"ad",  x"1a",  x"d0",  x"31", -- 1028
         x"d0",  x"d1",  x"e1",  x"a7",  x"ed",  x"52",  x"c3",  x"1a", -- 1030
         x"c9",  x"81",  x"bd",  x"2b",  x"d0",  x"d8",  x"cd",  x"2f", -- 1038
         x"d0",  x"74",  x"cc",  x"18",  x"cc",  x"81",  x"bc",  x"39", -- 1040
         x"d0",  x"4b",  x"d0",  x"d1",  x"e1",  x"7a",  x"ac",  x"17", -- 1048
         x"38",  x"03",  x"a7",  x"ed",  x"52",  x"cb",  x"7c",  x"20", -- 1050
         x"05",  x"21",  x"00",  x"00",  x"18",  x"03",  x"21",  x"01", -- 1058
         x"00",  x"c3",  x"1a",  x"c9",  x"82",  x"55",  x"bc",  x"45", -- 1060
         x"d0",  x"6b",  x"d0",  x"d1",  x"e1",  x"ed",  x"52",  x"21", -- 1068
         x"00",  x"00",  x"30",  x"01",  x"23",  x"c3",  x"1a",  x"c9", -- 1070
         x"81",  x"be",  x"64",  x"d0",  x"d8",  x"cd",  x"16",  x"cd", -- 1078
         x"49",  x"d0",  x"18",  x"cc",  x"83",  x"52",  x"4f",  x"d4", -- 1080
         x"78",  x"d0",  x"8c",  x"d0",  x"d1",  x"e1",  x"e3",  x"c3", -- 1088
         x"19",  x"c9",  x"85",  x"53",  x"50",  x"41",  x"43",  x"c5", -- 1090
         x"84",  x"d0",  x"d8",  x"cd",  x"77",  x"ce",  x"a5",  x"ca", -- 1098
         x"18",  x"cc",  x"84",  x"2d",  x"44",  x"55",  x"d0",  x"92", -- 10A0
         x"d0",  x"d8",  x"cd",  x"23",  x"cd",  x"68",  x"c9",  x"04", -- 10A8
         x"00",  x"23",  x"cd",  x"18",  x"cc",  x"88",  x"54",  x"52", -- 10B0
         x"41",  x"56",  x"45",  x"52",  x"53",  x"c5",  x"a2",  x"d0", -- 10B8
         x"d8",  x"cd",  x"16",  x"cd",  x"fa",  x"cc",  x"98",  x"cc", -- 10C0
         x"2c",  x"c9",  x"7f",  x"00",  x"fa",  x"cc",  x"73",  x"cd", -- 10C8
         x"49",  x"d0",  x"68",  x"c9",  x"f0",  x"ff",  x"16",  x"cd", -- 10D0
         x"09",  x"cd",  x"18",  x"cc",  x"86",  x"4c",  x"41",  x"54", -- 10D8
         x"45",  x"53",  x"d4",  x"b5",  x"d0",  x"d8",  x"cd",  x"7b", -- 10E0
         x"cf",  x"64",  x"cd",  x"64",  x"cd",  x"18",  x"cc",  x"83", -- 10E8
         x"4c",  x"46",  x"c1",  x"dc",  x"d0",  x"d8",  x"cd",  x"2c", -- 10F0
         x"c9",  x"04",  x"00",  x"2f",  x"d0",  x"18",  x"cc",  x"83", -- 10F8
         x"43",  x"46",  x"c1",  x"ef",  x"d0",  x"d8",  x"cd",  x"66", -- 1100
         x"ce",  x"2f",  x"d0",  x"18",  x"cc",  x"83",  x"4e",  x"46", -- 1108
         x"c1",  x"ff",  x"d0",  x"d8",  x"cd",  x"2c",  x"c9",  x"05", -- 1110
         x"00",  x"2f",  x"d0",  x"2c",  x"c9",  x"ff",  x"ff",  x"c0", -- 1118
         x"d0",  x"18",  x"cc",  x"83",  x"50",  x"46",  x"c1",  x"0d", -- 1120
         x"d1",  x"d8",  x"cd",  x"5e",  x"ce",  x"c0",  x"d0",  x"2c", -- 1128
         x"c9",  x"05",  x"00",  x"98",  x"cc",  x"18",  x"cc",  x"84", -- 1130
         x"21",  x"43",  x"53",  x"d0",  x"23",  x"d1",  x"d8",  x"cd", -- 1138
         x"ce",  x"cb",  x"b0",  x"cf",  x"95",  x"cd",  x"18",  x"cc", -- 1140
         x"86",  x"3f",  x"45",  x"52",  x"52",  x"4f",  x"d2",  x"37", -- 1148
         x"d1",  x"d8",  x"cd",  x"16",  x"cd",  x"68",  x"c9",  x"08", -- 1150
         x"00",  x"4c",  x"d6",  x"50",  x"c9",  x"04",  x"00",  x"09", -- 1158
         x"cd",  x"18",  x"cc",  x"85",  x"3f",  x"43",  x"4f",  x"4d", -- 1160
         x"d0",  x"48",  x"d1",  x"d8",  x"cd",  x"87",  x"cf",  x"64", -- 1168
         x"cd",  x"74",  x"cc",  x"2c",  x"c9",  x"11",  x"00",  x"51", -- 1170
         x"d1",  x"18",  x"cc",  x"85",  x"3f",  x"45",  x"58",  x"45", -- 1178
         x"c3",  x"63",  x"d1",  x"d8",  x"cd",  x"87",  x"cf",  x"64", -- 1180
         x"cd",  x"2c",  x"c9",  x"12",  x"00",  x"51",  x"d1",  x"18", -- 1188
         x"cc",  x"86",  x"3f",  x"50",  x"41",  x"49",  x"52",  x"d3", -- 1190
         x"7b",  x"d1",  x"d8",  x"cd",  x"2f",  x"d0",  x"2c",  x"c9", -- 1198
         x"13",  x"00",  x"51",  x"d1",  x"18",  x"cc",  x"84",  x"3f", -- 11A0
         x"43",  x"53",  x"d0",  x"91",  x"d1",  x"d8",  x"cd",  x"ce", -- 11A8
         x"cb",  x"b0",  x"cf",  x"64",  x"cd",  x"2f",  x"d0",  x"2c", -- 11B0
         x"c9",  x"14",  x"00",  x"51",  x"d1",  x"18",  x"cc",  x"88", -- 11B8
         x"3f",  x"4c",  x"4f",  x"41",  x"44",  x"49",  x"4e",  x"c7", -- 11C0
         x"a6",  x"d1",  x"d8",  x"cd",  x"42",  x"cf",  x"64",  x"cd", -- 11C8
         x"74",  x"cc",  x"2c",  x"c9",  x"16",  x"00",  x"51",  x"d1", -- 11D0
         x"18",  x"cc",  x"87",  x"43",  x"4f",  x"4d",  x"50",  x"49", -- 11D8
         x"4c",  x"c5",  x"bf",  x"d1",  x"d8",  x"cd",  x"6b",  x"d1", -- 11E0
         x"5a",  x"cc",  x"23",  x"cd",  x"e3",  x"cf",  x"45",  x"cc", -- 11E8
         x"64",  x"cd",  x"0e",  x"d0",  x"18",  x"cc",  x"c2",  x"28", -- 11F0
         x"a8",  x"da",  x"d1",  x"d8",  x"cd",  x"56",  x"ce",  x"87", -- 11F8
         x"cf",  x"95",  x"cd",  x"18",  x"cc",  x"82",  x"29",  x"a9", -- 1200
         x"f6",  x"d1",  x"d8",  x"cd",  x"2c",  x"c9",  x"c0",  x"00", -- 1208
         x"87",  x"cf",  x"95",  x"cd",  x"18",  x"cc",  x"86",  x"53", -- 1210
         x"4d",  x"55",  x"44",  x"47",  x"c5",  x"05",  x"d2",  x"d8", -- 1218
         x"cd",  x"e5",  x"d0",  x"2c",  x"c9",  x"20",  x"00",  x"56", -- 1220
         x"cd",  x"18",  x"cc",  x"83",  x"48",  x"45",  x"d8",  x"16", -- 1228
         x"d2",  x"d8",  x"cd",  x"2c",  x"c9",  x"10",  x"00",  x"92", -- 1230
         x"cf",  x"95",  x"cd",  x"18",  x"cc",  x"87",  x"44",  x"45", -- 1238
         x"43",  x"49",  x"4d",  x"41",  x"cc",  x"2b",  x"d2",  x"d8", -- 1240
         x"cd",  x"2c",  x"c9",  x"0a",  x"00",  x"92",  x"cf",  x"95", -- 1248
         x"cd",  x"18",  x"cc",  x"87",  x"28",  x"3b",  x"43",  x"4f", -- 1250
         x"44",  x"45",  x"a9",  x"3d",  x"d2",  x"d8",  x"cd",  x"5a", -- 1258
         x"cc",  x"e5",  x"d0",  x"29",  x"d1",  x"05",  x"d1",  x"95", -- 1260
         x"cd",  x"18",  x"cc",  x"c5",  x"3b",  x"43",  x"4f",  x"44", -- 1268
         x"c5",  x"53",  x"d2",  x"d8",  x"cd",  x"ad",  x"d1",  x"e4", -- 1270
         x"d1",  x"5d",  x"d2",  x"fb",  x"d1",  x"18",  x"cc",  x"87", -- 1278
         x"3c",  x"42",  x"55",  x"49",  x"4c",  x"44",  x"d3",  x"6b", -- 1280
         x"d2",  x"d8",  x"cd",  x"56",  x"ce",  x"05",  x"ce",  x"18", -- 1288
         x"cc",  x"85",  x"44",  x"4f",  x"45",  x"53",  x"be",  x"7f", -- 1290
         x"d2",  x"d8",  x"cd",  x"5a",  x"cc",  x"e5",  x"d0",  x"29", -- 1298
         x"d1",  x"95",  x"cd",  x"5d",  x"d2",  x"fd",  x"2b",  x"fd", -- 12A0
         x"70",  x"00",  x"fd",  x"2b",  x"fd",  x"71",  x"00",  x"13", -- 12A8
         x"eb",  x"4e",  x"23",  x"46",  x"23",  x"c3",  x"1a",  x"c9", -- 12B0
         x"85",  x"43",  x"4f",  x"55",  x"4e",  x"d4",  x"91",  x"d2", -- 12B8
         x"d8",  x"cd",  x"23",  x"cd",  x"d6",  x"cf",  x"16",  x"cd", -- 12C0
         x"73",  x"cd",  x"18",  x"cc",  x"84",  x"54",  x"59",  x"50", -- 12C8
         x"c5",  x"b8",  x"d2",  x"d8",  x"cd",  x"a9",  x"d0",  x"68", -- 12D0
         x"c9",  x"18",  x"00",  x"fa",  x"cc",  x"98",  x"cc",  x"16", -- 12D8
         x"cd",  x"cb",  x"c9",  x"e7",  x"c9",  x"73",  x"cd",  x"a5", -- 12E0
         x"ca",  x"7d",  x"c9",  x"f8",  x"ff",  x"50",  x"c9",  x"04", -- 12E8
         x"00",  x"09",  x"cd",  x"18",  x"cc",  x"89",  x"2d",  x"54", -- 12F0
         x"52",  x"41",  x"49",  x"4c",  x"49",  x"4e",  x"c7",  x"cc", -- 12F8
         x"d2",  x"d8",  x"cd",  x"23",  x"cd",  x"56",  x"ce",  x"cb", -- 1300
         x"c9",  x"fa",  x"cc",  x"fa",  x"cc",  x"98",  x"cc",  x"5e", -- 1308
         x"ce",  x"2f",  x"d0",  x"73",  x"cd",  x"77",  x"ce",  x"2f", -- 1310
         x"d0",  x"68",  x"c9",  x"08",  x"00",  x"2f",  x"cc",  x"50", -- 1318
         x"c9",  x"06",  x"00",  x"5e",  x"ce",  x"2f",  x"d0",  x"7d", -- 1320
         x"c9",  x"e0",  x"ff",  x"18",  x"cc",  x"84",  x"28",  x"2e", -- 1328
         x"22",  x"a9",  x"f5",  x"d2",  x"d8",  x"cd",  x"6d",  x"cc", -- 1330
         x"c0",  x"d2",  x"23",  x"cd",  x"d6",  x"cf",  x"5a",  x"cc", -- 1338
         x"98",  x"cc",  x"45",  x"cc",  x"d3",  x"d2",  x"18",  x"cc", -- 1340
         x"c2",  x"2e",  x"a2",  x"2d",  x"d3",  x"d8",  x"cd",  x"2c", -- 1348
         x"c9",  x"22",  x"00",  x"87",  x"cf",  x"64",  x"cd",  x"68", -- 1350
         x"c9",  x"14",  x"00",  x"e4",  x"d1",  x"34",  x"d3",  x"2e", -- 1358
         x"d5",  x"f2",  x"cf",  x"73",  x"cd",  x"d6",  x"cf",  x"02", -- 1360
         x"d0",  x"50",  x"c9",  x"0a",  x"00",  x"2e",  x"d5",  x"f2", -- 1368
         x"cf",  x"c0",  x"d2",  x"d3",  x"d2",  x"18",  x"cc",  x"88", -- 1370
         x"28",  x"45",  x"58",  x"50",  x"45",  x"43",  x"54",  x"a9", -- 1378
         x"48",  x"d3",  x"84",  x"d3",  x"d9",  x"cd",  x"4a",  x"02", -- 1380
         x"cd",  x"03",  x"f0",  x"16",  x"fe",  x"0d",  x"28",  x"06", -- 1388
         x"cd",  x"03",  x"f0",  x"00",  x"18",  x"f2",  x"ed",  x"5b", -- 1390
         x"a0",  x"b7",  x"7a",  x"b3",  x"28",  x"18",  x"3e",  x"08", -- 1398
         x"cd",  x"03",  x"f0",  x"00",  x"ed",  x"5b",  x"a0",  x"b7", -- 13A0
         x"cd",  x"03",  x"f0",  x"32",  x"7e",  x"b7",  x"20",  x"e6", -- 13A8
         x"3e",  x"09",  x"cd",  x"03",  x"f0",  x"00",  x"c1",  x"ed", -- 13B0
         x"5b",  x"a0",  x"b7",  x"cd",  x"03",  x"f0",  x"32",  x"56", -- 13B8
         x"78",  x"b1",  x"28",  x"11",  x"7a",  x"b7",  x"28",  x"0d", -- 13C0
         x"e1",  x"72",  x"23",  x"e5",  x"3e",  x"09",  x"cd",  x"03", -- 13C8
         x"f0",  x"00",  x"0b",  x"18",  x"e2",  x"3e",  x"09",  x"cd", -- 13D0
         x"03",  x"f0",  x"00",  x"e1",  x"36",  x"00",  x"cd",  x"51", -- 13D8
         x"02",  x"d9",  x"c3",  x"1b",  x"c9",  x"86",  x"45",  x"58", -- 13E0
         x"50",  x"45",  x"43",  x"d4",  x"77",  x"d3",  x"d8",  x"cd", -- 13E8
         x"2b",  x"cf",  x"73",  x"cd",  x"68",  x"c9",  x"6c",  x"00", -- 13F0
         x"fa",  x"cc",  x"98",  x"cc",  x"fa",  x"cc",  x"cb",  x"c9", -- 13F8
         x"c9",  x"ca",  x"23",  x"cd",  x"2c",  x"c9",  x"0e",  x"00", -- 1400
         x"a7",  x"ce",  x"64",  x"cd",  x"3d",  x"d0",  x"68",  x"c9", -- 1408
         x"20",  x"00",  x"09",  x"cd",  x"2c",  x"c9",  x"08",  x"00", -- 1410
         x"fa",  x"cc",  x"e7",  x"c9",  x"3d",  x"d0",  x"23",  x"cd", -- 1418
         x"5a",  x"cc",  x"66",  x"ce",  x"2f",  x"d0",  x"98",  x"cc", -- 1420
         x"45",  x"cc",  x"2f",  x"d0",  x"50",  x"c9",  x"28",  x"00", -- 1428
         x"23",  x"cd",  x"2c",  x"c9",  x"0d",  x"00",  x"3d",  x"d0", -- 1430
         x"68",  x"c9",  x"0e",  x"00",  x"2f",  x"cc",  x"09",  x"cd", -- 1438
         x"77",  x"ce",  x"56",  x"ce",  x"50",  x"c9",  x"04",  x"00", -- 1440
         x"23",  x"cd",  x"e7",  x"c9",  x"a4",  x"cd",  x"56",  x"ce", -- 1448
         x"e7",  x"c9",  x"d6",  x"cf",  x"95",  x"cd",  x"a5",  x"ca", -- 1450
         x"7d",  x"c9",  x"a6",  x"ff",  x"09",  x"cd",  x"50",  x"c9", -- 1458
         x"04",  x"00",  x"82",  x"d3",  x"18",  x"cc",  x"85",  x"51", -- 1460
         x"55",  x"45",  x"52",  x"d9",  x"e5",  x"d3",  x"d8",  x"cd", -- 1468
         x"c9",  x"ce",  x"64",  x"cd",  x"2c",  x"c9",  x"50",  x"00", -- 1470
         x"ee",  x"d3",  x"56",  x"ce",  x"4b",  x"cf",  x"95",  x"cd", -- 1478
         x"18",  x"cc",  x"c1",  x"80",  x"66",  x"d4",  x"d8",  x"cd", -- 1480
         x"42",  x"cf",  x"64",  x"cd",  x"68",  x"c9",  x"2a",  x"00", -- 1488
         x"5e",  x"ce",  x"42",  x"cf",  x"3f",  x"cd",  x"56",  x"ce", -- 1490
         x"4b",  x"cf",  x"95",  x"cd",  x"42",  x"cf",  x"64",  x"cd", -- 1498
         x"99",  x"ce",  x"5e",  x"ce",  x"2f",  x"d0",  x"96",  x"cb", -- 14A0
         x"74",  x"cc",  x"68",  x"c9",  x"08",  x"00",  x"83",  x"d1", -- 14A8
         x"5a",  x"cc",  x"09",  x"cd",  x"50",  x"c9",  x"06",  x"00", -- 14B0
         x"5a",  x"cc",  x"09",  x"cd",  x"18",  x"cc",  x"84",  x"46", -- 14B8
         x"49",  x"4c",  x"cc",  x"82",  x"d4",  x"c7",  x"d4",  x"69", -- 14C0
         x"60",  x"d1",  x"c1",  x"e3",  x"eb",  x"78",  x"b1",  x"28", -- 14C8
         x"06",  x"7d",  x"12",  x"13",  x"0b",  x"18",  x"f6",  x"c1", -- 14D0
         x"c3",  x"1b",  x"c9",  x"85",  x"45",  x"52",  x"41",  x"53", -- 14D8
         x"c5",  x"be",  x"d4",  x"d8",  x"cd",  x"56",  x"ce",  x"c5", -- 14E0
         x"d4",  x"18",  x"cc",  x"86",  x"42",  x"4c",  x"41",  x"4e", -- 14E8
         x"4b",  x"d3",  x"db",  x"d4",  x"d8",  x"cd",  x"77",  x"ce", -- 14F0
         x"c5",  x"d4",  x"18",  x"cc",  x"84",  x"48",  x"4f",  x"4c", -- 14F8
         x"c4",  x"eb",  x"d4",  x"d8",  x"cd",  x"2c",  x"c9",  x"ff", -- 1500
         x"ff",  x"c3",  x"cf",  x"3f",  x"cd",  x"c3",  x"cf",  x"64", -- 1508
         x"cd",  x"a4",  x"cd",  x"18",  x"cc",  x"83",  x"50",  x"41", -- 1510
         x"c4",  x"fc",  x"d4",  x"d8",  x"cd",  x"f2",  x"cf",  x"2c", -- 1518
         x"c9",  x"44",  x"00",  x"98",  x"cc",  x"18",  x"cc",  x"84", -- 1520
         x"57",  x"4f",  x"52",  x"c4",  x"15",  x"d5",  x"d8",  x"cd", -- 1528
         x"42",  x"cf",  x"64",  x"cd",  x"68",  x"c9",  x"0c",  x"00", -- 1530
         x"42",  x"cf",  x"64",  x"cd",  x"77",  x"db",  x"50",  x"c9", -- 1538
         x"06",  x"00",  x"c9",  x"ce",  x"64",  x"cd",  x"4b",  x"cf", -- 1540
         x"64",  x"cd",  x"98",  x"cc",  x"16",  x"cd",  x"6d",  x"ca", -- 1548
         x"f2",  x"cf",  x"2c",  x"c9",  x"22",  x"00",  x"f4",  x"d4", -- 1550
         x"4b",  x"cf",  x"3f",  x"cd",  x"fa",  x"cc",  x"2f",  x"d0", -- 1558
         x"45",  x"cc",  x"6d",  x"cc",  x"f2",  x"cf",  x"a4",  x"cd", -- 1560
         x"98",  x"cc",  x"f2",  x"cf",  x"d6",  x"cf",  x"5a",  x"cc", -- 1568
         x"13",  x"cb",  x"18",  x"cc",  x"88",  x"28",  x"4e",  x"55", -- 1570
         x"4d",  x"42",  x"45",  x"52",  x"a9",  x"27",  x"d5",  x"d8", -- 1578
         x"cd",  x"d6",  x"cf",  x"23",  x"cd",  x"45",  x"cc",  x"73", -- 1580
         x"cd",  x"92",  x"cf",  x"64",  x"cd",  x"fa",  x"c9",  x"68", -- 1588
         x"c9",  x"2c",  x"00",  x"16",  x"cd",  x"92",  x"cf",  x"64", -- 1590
         x"cd",  x"28",  x"cb",  x"09",  x"cd",  x"8a",  x"d0",  x"92", -- 1598
         x"cf",  x"64",  x"cd",  x"28",  x"cb",  x"a5",  x"cc",  x"9c", -- 15A0
         x"cf",  x"64",  x"cd",  x"d6",  x"cf",  x"68",  x"c9",  x"08", -- 15A8
         x"00",  x"5e",  x"ce",  x"9c",  x"cf",  x"3f",  x"cd",  x"5a", -- 15B0
         x"cc",  x"50",  x"c9",  x"c6",  x"ff",  x"5a",  x"cc",  x"18", -- 15B8
         x"cc",  x"86",  x"4e",  x"55",  x"4d",  x"42",  x"45",  x"d2", -- 15C0
         x"74",  x"d5",  x"d8",  x"cd",  x"56",  x"ce",  x"56",  x"ce", -- 15C8
         x"8a",  x"d0",  x"23",  x"cd",  x"d6",  x"cf",  x"73",  x"cd", -- 15D0
         x"2c",  x"c9",  x"2d",  x"00",  x"3d",  x"d0",  x"23",  x"cd", -- 15D8
         x"45",  x"cc",  x"98",  x"cc",  x"2c",  x"c9",  x"ff",  x"ff", -- 15E0
         x"9c",  x"cf",  x"95",  x"cd",  x"7f",  x"d5",  x"23",  x"cd", -- 15E8
         x"73",  x"cd",  x"77",  x"ce",  x"2f",  x"d0",  x"68",  x"c9", -- 15F0
         x"16",  x"00",  x"23",  x"cd",  x"73",  x"cd",  x"2c",  x"c9", -- 15F8
         x"2e",  x"00",  x"2f",  x"d0",  x"56",  x"ce",  x"51",  x"d1", -- 1600
         x"56",  x"ce",  x"50",  x"c9",  x"dc",  x"ff",  x"09",  x"cd", -- 1608
         x"5a",  x"cc",  x"68",  x"c9",  x"04",  x"00",  x"dd",  x"cc", -- 1610
         x"18",  x"cc",  x"85",  x"2d",  x"46",  x"49",  x"4e",  x"c4", -- 1618
         x"c1",  x"d5",  x"d8",  x"cd",  x"77",  x"ce",  x"2e",  x"d5", -- 1620
         x"f2",  x"cf",  x"6d",  x"cf",  x"64",  x"cd",  x"64",  x"cd", -- 1628
         x"23",  x"ca",  x"23",  x"cd",  x"74",  x"cc",  x"68",  x"c9", -- 1630
         x"0a",  x"00",  x"09",  x"cd",  x"f2",  x"cf",  x"e5",  x"d0", -- 1638
         x"23",  x"ca",  x"18",  x"cc",  x"85",  x"45",  x"52",  x"52", -- 1640
         x"4f",  x"d2",  x"1a",  x"d6",  x"d8",  x"cd",  x"e3",  x"ce", -- 1648
         x"64",  x"cd",  x"87",  x"cc",  x"68",  x"c9",  x"04",  x"00", -- 1650
         x"62",  x"02",  x"f2",  x"cf",  x"c0",  x"d2",  x"d3",  x"d2", -- 1658
         x"34",  x"d3",  x"02",  x"3f",  x"20",  x"c7",  x"da",  x"dd", -- 1660
         x"cb",  x"42",  x"cf",  x"64",  x"cd",  x"a9",  x"d0",  x"68", -- 1668
         x"c9",  x"08",  x"00",  x"4b",  x"cf",  x"64",  x"cd",  x"16", -- 1670
         x"cd",  x"52",  x"d8",  x"83",  x"49",  x"44",  x"ae",  x"44", -- 1678
         x"d6",  x"d8",  x"cd",  x"1b",  x"d5",  x"2c",  x"c9",  x"20", -- 1680
         x"00",  x"2c",  x"c9",  x"5f",  x"00",  x"c5",  x"d4",  x"23", -- 1688
         x"cd",  x"29",  x"d1",  x"f5",  x"d0",  x"fa",  x"cc",  x"2f", -- 1690
         x"d0",  x"1b",  x"d5",  x"16",  x"cd",  x"13",  x"cb",  x"1b", -- 1698
         x"d5",  x"c0",  x"d2",  x"2c",  x"c9",  x"1f",  x"00",  x"96", -- 16A0
         x"cb",  x"d3",  x"d2",  x"9a",  x"d0",  x"18",  x"cc",  x"86", -- 16A8
         x"43",  x"52",  x"45",  x"41",  x"54",  x"c5",  x"7b",  x"d6", -- 16B0
         x"d8",  x"cd",  x"22",  x"d6",  x"68",  x"c9",  x"10",  x"00", -- 16B8
         x"09",  x"cd",  x"13",  x"d1",  x"81",  x"d6",  x"2c",  x"c9", -- 16C0
         x"04",  x"00",  x"c7",  x"da",  x"9a",  x"d0",  x"f2",  x"cf", -- 16C8
         x"23",  x"cd",  x"73",  x"cd",  x"d5",  x"ce",  x"64",  x"cd", -- 16D0
         x"96",  x"d9",  x"d6",  x"cf",  x"02",  x"d0",  x"23",  x"cd", -- 16D8
         x"2c",  x"c9",  x"a0",  x"00",  x"56",  x"cd",  x"f2",  x"cf", -- 16E0
         x"5e",  x"ce",  x"2f",  x"d0",  x"2c",  x"c9",  x"80",  x"00", -- 16E8
         x"56",  x"cd",  x"e5",  x"d0",  x"0e",  x"d0",  x"7b",  x"cf", -- 16F0
         x"64",  x"cd",  x"95",  x"cd",  x"f2",  x"cf",  x"e3",  x"cf", -- 16F8
         x"0e",  x"d0",  x"18",  x"cc",  x"c9",  x"28",  x"43",  x"4f", -- 1700
         x"4d",  x"50",  x"49",  x"4c",  x"45",  x"a9",  x"af",  x"d6", -- 1708
         x"d8",  x"cd",  x"22",  x"d6",  x"74",  x"cc",  x"56",  x"ce", -- 1710
         x"51",  x"d1",  x"09",  x"cd",  x"05",  x"d1",  x"0e",  x"d0", -- 1718
         x"18",  x"cc",  x"c7",  x"4c",  x"49",  x"54",  x"45",  x"52", -- 1720
         x"41",  x"cc",  x"04",  x"d7",  x"d8",  x"cd",  x"87",  x"cf", -- 1728
         x"64",  x"cd",  x"68",  x"c9",  x"08",  x"00",  x"e4",  x"d1", -- 1730
         x"2c",  x"c9",  x"0e",  x"d0",  x"18",  x"cc",  x"c8",  x"44", -- 1738
         x"4c",  x"49",  x"54",  x"45",  x"52",  x"41",  x"cc",  x"22", -- 1740
         x"d7",  x"d8",  x"cd",  x"87",  x"cf",  x"64",  x"cd",  x"68", -- 1748
         x"c9",  x"08",  x"00",  x"16",  x"cd",  x"2c",  x"d7",  x"2c", -- 1750
         x"d7",  x"18",  x"cc",  x"86",  x"3f",  x"53",  x"54",  x"41", -- 1758
         x"43",  x"cb",  x"3e",  x"d7",  x"d8",  x"cd",  x"ce",  x"cb", -- 1760
         x"b6",  x"ce",  x"64",  x"cd",  x"16",  x"cd",  x"69",  x"d0", -- 1768
         x"5e",  x"ce",  x"51",  x"d1",  x"ce",  x"cb",  x"56",  x"ce", -- 1770
         x"2c",  x"c9",  x"20",  x"00",  x"98",  x"cc",  x"69",  x"d0", -- 1778
         x"2c",  x"c9",  x"07",  x"00",  x"51",  x"d1",  x"18",  x"cc", -- 1780
         x"89",  x"49",  x"4e",  x"54",  x"45",  x"52",  x"50",  x"52", -- 1788
         x"45",  x"d4",  x"5b",  x"d7",  x"d8",  x"cd",  x"22",  x"d6", -- 1790
         x"68",  x"c9",  x"1e",  x"00",  x"87",  x"cf",  x"64",  x"cd", -- 1798
         x"49",  x"d0",  x"68",  x"c9",  x"0a",  x"00",  x"05",  x"d1", -- 17A0
         x"0e",  x"d0",  x"50",  x"c9",  x"06",  x"00",  x"05",  x"d1", -- 17A8
         x"41",  x"c9",  x"64",  x"d7",  x"50",  x"c9",  x"1c",  x"00", -- 17B0
         x"f2",  x"cf",  x"ca",  x"d5",  x"9c",  x"cf",  x"64",  x"cd", -- 17B8
         x"d6",  x"cf",  x"68",  x"c9",  x"08",  x"00",  x"49",  x"d7", -- 17C0
         x"50",  x"c9",  x"06",  x"00",  x"09",  x"cd",  x"2c",  x"d7", -- 17C8
         x"64",  x"d7",  x"50",  x"c9",  x"c2",  x"ff",  x"89",  x"49", -- 17D0
         x"4d",  x"4d",  x"45",  x"44",  x"49",  x"41",  x"54",  x"c5", -- 17D8
         x"88",  x"d7",  x"d8",  x"cd",  x"e5",  x"d0",  x"2c",  x"c9", -- 17E0
         x"40",  x"00",  x"56",  x"cd",  x"18",  x"cc",  x"8a",  x"56", -- 17E8
         x"4f",  x"43",  x"41",  x"42",  x"55",  x"4c",  x"41",  x"52", -- 17F0
         x"d9",  x"d6",  x"d7",  x"d8",  x"cd",  x"89",  x"d2",  x"2c", -- 17F8
         x"c9",  x"81",  x"a0",  x"0e",  x"d0",  x"7b",  x"cf",  x"64", -- 1800
         x"cd",  x"05",  x"d1",  x"0e",  x"d0",  x"f2",  x"cf",  x"07", -- 1808
         x"cf",  x"64",  x"cd",  x"0e",  x"d0",  x"07",  x"cf",  x"95", -- 1810
         x"cd",  x"99",  x"d2",  x"e3",  x"cf",  x"6d",  x"cf",  x"95", -- 1818
         x"cd",  x"18",  x"cc",  x"8b",  x"44",  x"45",  x"46",  x"49", -- 1820
         x"4e",  x"49",  x"54",  x"49",  x"4f",  x"4e",  x"d3",  x"ee", -- 1828
         x"d7",  x"d8",  x"cd",  x"6d",  x"cf",  x"64",  x"cd",  x"7b", -- 1830
         x"cf",  x"95",  x"cd",  x"18",  x"cc",  x"c1",  x"a8",  x"23", -- 1838
         x"d8",  x"d8",  x"cd",  x"2c",  x"c9",  x"29",  x"00",  x"2e", -- 1840
         x"d5",  x"18",  x"cc",  x"84",  x"51",  x"55",  x"49",  x"d4", -- 1848
         x"3d",  x"d8",  x"d8",  x"cd",  x"56",  x"ce",  x"42",  x"cf", -- 1850
         x"95",  x"cd",  x"fb",  x"d1",  x"01",  x"cc",  x"fa",  x"ca", -- 1858
         x"6e",  x"d4",  x"94",  x"d7",  x"87",  x"cf",  x"64",  x"cd", -- 1860
         x"74",  x"cc",  x"68",  x"c9",  x"07",  x"00",  x"34",  x"d3", -- 1868
         x"02",  x"4f",  x"4b",  x"50",  x"c9",  x"e7",  x"ff",  x"85", -- 1870
         x"41",  x"42",  x"4f",  x"52",  x"d4",  x"4b",  x"d8",  x"d8", -- 1878
         x"cd",  x"dd",  x"cb",  x"47",  x"d2",  x"64",  x"d7",  x"fa", -- 1880
         x"ca",  x"34",  x"d3",  x"0e",  x"4b",  x"43",  x"20",  x"2d", -- 1888
         x"20",  x"46",  x"4f",  x"52",  x"54",  x"48",  x"20",  x"33", -- 1890
         x"2e",  x"31",  x"70",  x"02",  x"31",  x"d8",  x"52",  x"d8", -- 1898
         x"84",  x"57",  x"41",  x"52",  x"cd",  x"77",  x"d8",  x"d8", -- 18A0
         x"cd",  x"4f",  x"db",  x"7f",  x"d8",  x"84",  x"43",  x"4f", -- 18A8
         x"4c",  x"c4",  x"a0",  x"d8",  x"cc",  x"d8",  x"01",  x"ca", -- 18B0
         x"d8",  x"2a",  x"2a",  x"c0",  x"f9",  x"2a",  x"28",  x"c0", -- 18B8
         x"22",  x"7e",  x"01",  x"fd",  x"2a",  x"2c",  x"c0",  x"c3", -- 18C0
         x"1b",  x"c9",  x"a7",  x"d8",  x"21",  x"f7",  x"d8",  x"11", -- 18C8
         x"4a",  x"02",  x"01",  x"43",  x"00",  x"ed",  x"b0",  x"2a", -- 18D0
         x"28",  x"c0",  x"11",  x"06",  x"00",  x"19",  x"54",  x"5d", -- 18D8
         x"21",  x"2a",  x"c0",  x"01",  x"18",  x"00",  x"ed",  x"b0", -- 18E0
         x"2a",  x"bb",  x"b7",  x"22",  x"48",  x"02",  x"1e",  x"24", -- 18E8
         x"3e",  x"0c",  x"cd",  x"0c",  x"f0",  x"18",  x"bf",  x"db", -- 18F0
         x"88",  x"cb",  x"d7",  x"d3",  x"88",  x"c9",  x"db",  x"88", -- 18F8
         x"cb",  x"97",  x"d3",  x"88",  x"c9",  x"87",  x"28",  x"41", -- 1900
         x"42",  x"4f",  x"52",  x"54",  x"a9",  x"ad",  x"d8",  x"d8", -- 1908
         x"cd",  x"7f",  x"d8",  x"18",  x"cc",  x"c5",  x"46",  x"4f", -- 1910
         x"52",  x"54",  x"c8",  x"58",  x"02",  x"a5",  x"d2",  x"1b", -- 1918
         x"d8",  x"81",  x"a0",  x"10",  x"c9",  x"00",  x"00",  x"c6", -- 1920
         x"45",  x"44",  x"49",  x"54",  x"4f",  x"d2",  x"68",  x"02", -- 1928
         x"a5",  x"d2",  x"1b",  x"d8",  x"81",  x"a0",  x"a3",  x"c7", -- 1930
         x"78",  x"02",  x"84",  x"53",  x"2d",  x"3e",  x"c4",  x"7a", -- 1938
         x"02",  x"43",  x"d9",  x"d1",  x"21",  x"00",  x"00",  x"7a", -- 1940
         x"e6",  x"80",  x"28",  x"01",  x"2b",  x"c3",  x"19",  x"c9", -- 1948
         x"82",  x"2b",  x"ad",  x"3a",  x"d9",  x"d8",  x"cd",  x"87", -- 1950
         x"cc",  x"68",  x"c9",  x"04",  x"00",  x"c8",  x"cc",  x"18", -- 1958
         x"cc",  x"83",  x"44",  x"2b",  x"ad",  x"50",  x"d9",  x"d8", -- 1960
         x"cd",  x"87",  x"cc",  x"68",  x"c9",  x"04",  x"00",  x"dd", -- 1968
         x"cc",  x"18",  x"cc",  x"83",  x"41",  x"42",  x"d3",  x"61", -- 1970
         x"d9",  x"d8",  x"cd",  x"23",  x"cd",  x"55",  x"d9",  x"18", -- 1978
         x"cc",  x"84",  x"44",  x"41",  x"42",  x"d3",  x"73",  x"d9", -- 1980
         x"d8",  x"cd",  x"23",  x"cd",  x"67",  x"d9",  x"18",  x"cc", -- 1988
         x"83",  x"4d",  x"49",  x"ce",  x"81",  x"d9",  x"d8",  x"cd", -- 1990
         x"31",  x"cd",  x"7c",  x"d0",  x"68",  x"c9",  x"04",  x"00", -- 1998
         x"16",  x"cd",  x"09",  x"cd",  x"18",  x"cc",  x"83",  x"4d", -- 19A0
         x"41",  x"d8",  x"90",  x"d9",  x"d8",  x"cd",  x"31",  x"cd", -- 19A8
         x"49",  x"d0",  x"68",  x"c9",  x"04",  x"00",  x"16",  x"cd", -- 19B0
         x"09",  x"cd",  x"18",  x"cc",  x"82",  x"4d",  x"aa",  x"a6", -- 19B8
         x"d9",  x"d8",  x"cd",  x"31",  x"cd",  x"bb",  x"cb",  x"45", -- 19C0
         x"cc",  x"79",  x"d9",  x"16",  x"cd",  x"79",  x"d9",  x"28", -- 19C8
         x"cb",  x"5a",  x"cc",  x"67",  x"d9",  x"18",  x"cc",  x"82", -- 19D0
         x"4d",  x"af",  x"bc",  x"d9",  x"d8",  x"cd",  x"fa",  x"cc", -- 19D8
         x"45",  x"cc",  x"45",  x"cc",  x"88",  x"d9",  x"6d",  x"cc", -- 19E0
         x"79",  x"d9",  x"54",  x"cb",  x"5a",  x"cc",  x"6d",  x"cc", -- 19E8
         x"bb",  x"cb",  x"55",  x"d9",  x"16",  x"cd",  x"5a",  x"cc", -- 19F0
         x"55",  x"d9",  x"16",  x"cd",  x"18",  x"cc",  x"81",  x"aa", -- 19F8
         x"d7",  x"d9",  x"d8",  x"cd",  x"c1",  x"d9",  x"09",  x"cd", -- 1A00
         x"18",  x"cc",  x"84",  x"2f",  x"4d",  x"4f",  x"c4",  x"fe", -- 1A08
         x"d9",  x"d8",  x"cd",  x"45",  x"cc",  x"41",  x"d9",  x"5a", -- 1A10
         x"cc",  x"dc",  x"d9",  x"18",  x"cc",  x"81",  x"af",  x"0a", -- 1A18
         x"da",  x"d8",  x"cd",  x"11",  x"da",  x"16",  x"cd",  x"09", -- 1A20
         x"cd",  x"18",  x"cc",  x"83",  x"4d",  x"4f",  x"c4",  x"1d", -- 1A28
         x"da",  x"d8",  x"cd",  x"11",  x"da",  x"09",  x"cd",  x"18", -- 1A30
         x"cc",  x"85",  x"2a",  x"2f",  x"4d",  x"4f",  x"c4",  x"2b", -- 1A38
         x"da",  x"d8",  x"cd",  x"45",  x"cc",  x"c1",  x"d9",  x"5a", -- 1A40
         x"cc",  x"dc",  x"d9",  x"18",  x"cc",  x"82",  x"2a",  x"af", -- 1A48
         x"39",  x"da",  x"d8",  x"cd",  x"41",  x"da",  x"16",  x"cd", -- 1A50
         x"09",  x"cd",  x"18",  x"cc",  x"85",  x"4d",  x"2f",  x"4d", -- 1A58
         x"4f",  x"c4",  x"4d",  x"da",  x"d8",  x"cd",  x"45",  x"cc", -- 1A60
         x"56",  x"ce",  x"6d",  x"cc",  x"54",  x"cb",  x"5a",  x"cc", -- 1A68
         x"16",  x"cd",  x"45",  x"cc",  x"54",  x"cb",  x"5a",  x"cc", -- 1A70
         x"18",  x"cc",  x"86",  x"28",  x"4c",  x"49",  x"4e",  x"45", -- 1A78
         x"a9",  x"5c",  x"da",  x"d8",  x"cd",  x"2c",  x"c9",  x"10", -- 1A80
         x"00",  x"02",  x"da",  x"98",  x"cc",  x"2c",  x"c9",  x"10", -- 1A88
         x"00",  x"11",  x"da",  x"45",  x"cc",  x"81",  x"ce",  x"8d", -- 1A90
         x"ce",  x"41",  x"da",  x"5a",  x"cc",  x"99",  x"ce",  x"02", -- 1A98
         x"da",  x"98",  x"cc",  x"77",  x"db",  x"98",  x"cc",  x"81", -- 1AA0
         x"ce",  x"18",  x"cc",  x"85",  x"2e",  x"4c",  x"49",  x"4e", -- 1AA8
         x"c5",  x"7a",  x"da",  x"d8",  x"cd",  x"83",  x"da",  x"01", -- 1AB0
         x"d3",  x"d3",  x"d2",  x"18",  x"cc",  x"87",  x"4d",  x"45", -- 1AB8
         x"53",  x"53",  x"41",  x"47",  x"c5",  x"ab",  x"da",  x"d8", -- 1AC0
         x"cd",  x"e3",  x"ce",  x"64",  x"cd",  x"68",  x"c9",  x"12", -- 1AC8
         x"00",  x"a9",  x"d0",  x"68",  x"c9",  x"08",  x"00",  x"5e", -- 1AD0
         x"ce",  x"b3",  x"da",  x"9a",  x"d0",  x"50",  x"c9",  x"0d", -- 1AD8
         x"00",  x"34",  x"d3",  x"06",  x"4d",  x"53",  x"47",  x"20", -- 1AE0
         x"23",  x"20",  x"5e",  x"de",  x"18",  x"cc",  x"87",  x"52", -- 1AE8
         x"45",  x"43",  x"2f",  x"42",  x"4c",  x"cb",  x"bd",  x"da", -- 1AF0
         x"0f",  x"ce",  x"04",  x"00",  x"85",  x"23",  x"42",  x"55", -- 1AF8
         x"46",  x"c6",  x"ee",  x"da",  x"d8",  x"cd",  x"1f",  x"cf", -- 1B00
         x"64",  x"cd",  x"13",  x"cf",  x"64",  x"cd",  x"2f",  x"d0", -- 1B08
         x"56",  x"ce",  x"8d",  x"ce",  x"e3",  x"cf",  x"54",  x"cb", -- 1B10
         x"16",  x"cd",  x"09",  x"cd",  x"18",  x"cc",  x"8d",  x"45", -- 1B18
         x"4d",  x"50",  x"54",  x"59",  x"2d",  x"42",  x"55",  x"46", -- 1B20
         x"46",  x"45",  x"52",  x"d3",  x"fc",  x"da",  x"d8",  x"cd", -- 1B28
         x"13",  x"cf",  x"64",  x"cd",  x"1f",  x"cf",  x"64",  x"cd", -- 1B30
         x"fa",  x"cc",  x"2f",  x"d0",  x"e3",  x"d4",  x"18",  x"cc", -- 1B38
         x"8c",  x"49",  x"4e",  x"49",  x"54",  x"2d",  x"42",  x"55", -- 1B40
         x"46",  x"46",  x"45",  x"52",  x"d3",  x"1e",  x"db",  x"d8", -- 1B48
         x"cd",  x"1f",  x"cf",  x"64",  x"cd",  x"13",  x"cf",  x"64", -- 1B50
         x"cd",  x"8d",  x"ce",  x"98",  x"cc",  x"cb",  x"c9",  x"56", -- 1B58
         x"ce",  x"e7",  x"c9",  x"95",  x"cd",  x"8d",  x"ce",  x"e3", -- 1B60
         x"cf",  x"bf",  x"c9",  x"f4",  x"ff",  x"18",  x"cc",  x"85", -- 1B68
         x"42",  x"4c",  x"4f",  x"43",  x"cb",  x"40",  x"db",  x"d8", -- 1B70
         x"cd",  x"5e",  x"ce",  x"ac",  x"d9",  x"04",  x"db",  x"96", -- 1B78
         x"d9",  x"5e",  x"ce",  x"2f",  x"d0",  x"8d",  x"ce",  x"e3", -- 1B80
         x"cf",  x"02",  x"da",  x"13",  x"cf",  x"64",  x"cd",  x"98", -- 1B88
         x"cc",  x"18",  x"cc",  x"84",  x"4c",  x"4f",  x"41",  x"c4", -- 1B90
         x"6f",  x"db",  x"d8",  x"cd",  x"42",  x"cf",  x"64",  x"cd", -- 1B98
         x"45",  x"cc",  x"4b",  x"cf",  x"64",  x"cd",  x"45",  x"cc", -- 1BA0
         x"56",  x"ce",  x"4b",  x"cf",  x"95",  x"cd",  x"99",  x"ce", -- 1BA8
         x"02",  x"da",  x"42",  x"cf",  x"95",  x"cd",  x"94",  x"d7", -- 1BB0
         x"5a",  x"cc",  x"4b",  x"cf",  x"95",  x"cd",  x"5a",  x"cc", -- 1BB8
         x"42",  x"cf",  x"95",  x"cd",  x"18",  x"cc",  x"c3",  x"2d", -- 1BC0
         x"2d",  x"be",  x"93",  x"db",  x"d8",  x"cd",  x"ca",  x"d1", -- 1BC8
         x"56",  x"ce",  x"4b",  x"cf",  x"95",  x"cd",  x"99",  x"ce", -- 1BD0
         x"42",  x"cf",  x"64",  x"cd",  x"fa",  x"cc",  x"31",  x"da", -- 1BD8
         x"2f",  x"d0",  x"42",  x"cf",  x"3f",  x"cd",  x"18",  x"cc", -- 1BE0
         x"c1",  x"a7",  x"c6",  x"db",  x"d8",  x"cd",  x"22",  x"d6", -- 1BE8
         x"74",  x"cc",  x"56",  x"ce",  x"51",  x"d1",  x"09",  x"cd", -- 1BF0
         x"2c",  x"d7",  x"18",  x"cc",  x"86",  x"46",  x"4f",  x"52", -- 1BF8
         x"47",  x"45",  x"d4",  x"e8",  x"db",  x"d8",  x"cd",  x"ec", -- 1C00
         x"db",  x"13",  x"d1",  x"23",  x"cd",  x"ef",  x"ce",  x"64", -- 1C08
         x"cd",  x"49",  x"d0",  x"2c",  x"c9",  x"15",  x"00",  x"51", -- 1C10
         x"d1",  x"45",  x"cc",  x"07",  x"cf",  x"64",  x"cd",  x"6d", -- 1C18
         x"cc",  x"fa",  x"cc",  x"49",  x"d0",  x"68",  x"c9",  x"12", -- 1C20
         x"00",  x"70",  x"02",  x"31",  x"d8",  x"64",  x"cd",  x"23", -- 1C28
         x"cd",  x"07",  x"cf",  x"95",  x"cd",  x"50",  x"c9",  x"e8", -- 1C30
         x"ff",  x"23",  x"cd",  x"2c",  x"c9",  x"04",  x"00",  x"2f", -- 1C38
         x"d0",  x"29",  x"d1",  x"f5",  x"d0",  x"64",  x"cd",  x"23", -- 1C40
         x"cd",  x"6d",  x"cc",  x"49",  x"d0",  x"68",  x"c9",  x"f2", -- 1C48
         x"ff",  x"fa",  x"cc",  x"66",  x"ce",  x"2f",  x"d0",  x"95", -- 1C50
         x"cd",  x"64",  x"cd",  x"a9",  x"d0",  x"74",  x"cc",  x"68", -- 1C58
         x"c9",  x"d8",  x"ff",  x"5a",  x"cc",  x"f8",  x"ce",  x"95", -- 1C60
         x"cd",  x"18",  x"cc",  x"84",  x"42",  x"41",  x"43",  x"cb", -- 1C68
         x"fc",  x"db",  x"d8",  x"cd",  x"f2",  x"cf",  x"2f",  x"d0", -- 1C70
         x"0e",  x"d0",  x"18",  x"cc",  x"c5",  x"42",  x"45",  x"47", -- 1C78
         x"49",  x"ce",  x"6b",  x"dc",  x"d8",  x"cd",  x"6b",  x"d1", -- 1C80
         x"f2",  x"cf",  x"5e",  x"ce",  x"18",  x"cc",  x"c5",  x"45", -- 1C88
         x"4e",  x"44",  x"49",  x"c6",  x"7c",  x"dc",  x"d8",  x"cd", -- 1C90
         x"6b",  x"d1",  x"66",  x"ce",  x"9a",  x"d1",  x"f2",  x"cf", -- 1C98
         x"fa",  x"cc",  x"2f",  x"d0",  x"16",  x"cd",  x"95",  x"cd", -- 1CA0
         x"18",  x"cc",  x"c2",  x"44",  x"cf",  x"8e",  x"dc",  x"d8", -- 1CA8
         x"cd",  x"e4",  x"d1",  x"cb",  x"c9",  x"f2",  x"cf",  x"6e", -- 1CB0
         x"ce",  x"18",  x"cc",  x"c4",  x"4c",  x"4f",  x"4f",  x"d0", -- 1CB8
         x"aa",  x"dc",  x"d8",  x"cd",  x"6e",  x"ce",  x"9a",  x"d1", -- 1CC0
         x"e4",  x"d1",  x"7d",  x"c9",  x"72",  x"dc",  x"18",  x"cc", -- 1CC8
         x"c5",  x"2b",  x"4c",  x"4f",  x"4f",  x"d0",  x"bb",  x"dc", -- 1CD0
         x"d8",  x"cd",  x"6e",  x"ce",  x"9a",  x"d1",  x"e4",  x"d1", -- 1CD8
         x"bf",  x"c9",  x"72",  x"dc",  x"18",  x"cc",  x"c5",  x"55", -- 1CE0
         x"4e",  x"54",  x"49",  x"cc",  x"d0",  x"dc",  x"d8",  x"cd", -- 1CE8
         x"5e",  x"ce",  x"9a",  x"d1",  x"e4",  x"d1",  x"68",  x"c9", -- 1CF0
         x"72",  x"dc",  x"18",  x"cc",  x"c5",  x"41",  x"47",  x"41", -- 1CF8
         x"49",  x"ce",  x"e6",  x"dc",  x"d8",  x"cd",  x"5e",  x"ce", -- 1D00
         x"9a",  x"d1",  x"e4",  x"d1",  x"50",  x"c9",  x"72",  x"dc", -- 1D08
         x"18",  x"cc",  x"c6",  x"52",  x"45",  x"50",  x"45",  x"41", -- 1D10
         x"d4",  x"fc",  x"dc",  x"d8",  x"cd",  x"45",  x"cc",  x"45", -- 1D18
         x"cc",  x"04",  x"dd",  x"5a",  x"cc",  x"5a",  x"cc",  x"66", -- 1D20
         x"ce",  x"2f",  x"d0",  x"96",  x"dc",  x"18",  x"cc",  x"c2", -- 1D28
         x"49",  x"c6",  x"12",  x"dd",  x"d8",  x"cd",  x"e4",  x"d1", -- 1D30
         x"68",  x"c9",  x"f2",  x"cf",  x"56",  x"ce",  x"0e",  x"d0", -- 1D38
         x"66",  x"ce",  x"18",  x"cc",  x"c4",  x"45",  x"4c",  x"53", -- 1D40
         x"c5",  x"2f",  x"dd",  x"d8",  x"cd",  x"66",  x"ce",  x"9a", -- 1D48
         x"d1",  x"e4",  x"d1",  x"50",  x"c9",  x"f2",  x"cf",  x"56", -- 1D50
         x"ce",  x"0e",  x"d0",  x"16",  x"cd",  x"66",  x"ce",  x"96", -- 1D58
         x"dc",  x"66",  x"ce",  x"18",  x"cc",  x"c5",  x"57",  x"48", -- 1D60
         x"49",  x"4c",  x"c5",  x"44",  x"dd",  x"d8",  x"cd",  x"34", -- 1D68
         x"dd",  x"e3",  x"cf",  x"18",  x"cc",  x"86",  x"53",  x"50", -- 1D70
         x"41",  x"43",  x"45",  x"d3",  x"65",  x"dd",  x"d8",  x"cd", -- 1D78
         x"56",  x"ce",  x"ac",  x"d9",  x"a9",  x"d0",  x"68",  x"c9", -- 1D80
         x"0c",  x"00",  x"56",  x"ce",  x"cb",  x"c9",  x"9a",  x"d0", -- 1D88
         x"7d",  x"c9",  x"fc",  x"ff",  x"18",  x"cc",  x"82",  x"3c", -- 1D90
         x"a3",  x"75",  x"dd",  x"d8",  x"cd",  x"1b",  x"d5",  x"c3", -- 1D98
         x"cf",  x"95",  x"cd",  x"18",  x"cc",  x"82",  x"23",  x"be", -- 1DA0
         x"96",  x"dd",  x"d8",  x"cd",  x"09",  x"cd",  x"09",  x"cd", -- 1DA8
         x"c3",  x"cf",  x"64",  x"cd",  x"1b",  x"d5",  x"fa",  x"cc", -- 1DB0
         x"2f",  x"d0",  x"18",  x"cc",  x"84",  x"53",  x"49",  x"47", -- 1DB8
         x"ce",  x"a5",  x"dd",  x"d8",  x"cd",  x"8a",  x"d0",  x"87", -- 1DC0
         x"cc",  x"68",  x"c9",  x"08",  x"00",  x"2c",  x"c9",  x"2d", -- 1DC8
         x"00",  x"03",  x"d5",  x"18",  x"cc",  x"81",  x"a3",  x"bc", -- 1DD0
         x"dd",  x"d8",  x"cd",  x"92",  x"cf",  x"64",  x"cd",  x"64", -- 1DD8
         x"da",  x"8a",  x"d0",  x"2c",  x"c9",  x"09",  x"00",  x"fa", -- 1DE0
         x"cc",  x"49",  x"d0",  x"68",  x"c9",  x"08",  x"00",  x"2c", -- 1DE8
         x"c9",  x"07",  x"00",  x"98",  x"cc",  x"2c",  x"c9",  x"30", -- 1DF0
         x"00",  x"98",  x"cc",  x"03",  x"d5",  x"18",  x"cc",  x"82", -- 1DF8
         x"23",  x"d3",  x"d5",  x"dd",  x"d8",  x"cd",  x"d9",  x"dd", -- 1E00
         x"fa",  x"cc",  x"fa",  x"cc",  x"a8",  x"cb",  x"74",  x"cc", -- 1E08
         x"68",  x"c9",  x"f4",  x"ff",  x"18",  x"cc",  x"83",  x"44", -- 1E10
         x"2e",  x"d2",  x"ff",  x"dd",  x"d8",  x"cd",  x"45",  x"cc", -- 1E18
         x"16",  x"cd",  x"fa",  x"cc",  x"88",  x"d9",  x"9b",  x"dd", -- 1E20
         x"04",  x"de",  x"c3",  x"dd",  x"aa",  x"dd",  x"5a",  x"cc", -- 1E28
         x"fa",  x"cc",  x"2f",  x"d0",  x"7e",  x"dd",  x"d3",  x"d2", -- 1E30
         x"18",  x"cc",  x"82",  x"2e",  x"d2",  x"16",  x"de",  x"d8", -- 1E38
         x"cd",  x"45",  x"cc",  x"41",  x"d9",  x"5a",  x"cc",  x"1c", -- 1E40
         x"de",  x"18",  x"cc",  x"82",  x"44",  x"ae",  x"3a",  x"de", -- 1E48
         x"d8",  x"cd",  x"56",  x"ce",  x"1c",  x"de",  x"9a",  x"d0", -- 1E50
         x"18",  x"cc",  x"81",  x"ae",  x"4b",  x"de",  x"d8",  x"cd", -- 1E58
         x"41",  x"d9",  x"50",  x"de",  x"18",  x"cc",  x"81",  x"bf", -- 1E60
         x"5a",  x"de",  x"d8",  x"cd",  x"64",  x"cd",  x"5e",  x"de", -- 1E68
         x"18",  x"cc",  x"82",  x"55",  x"ae",  x"66",  x"de",  x"d8", -- 1E70
         x"cd",  x"56",  x"ce",  x"50",  x"de",  x"18",  x"cc",  x"85", -- 1E78
         x"56",  x"4c",  x"49",  x"53",  x"d4",  x"72",  x"de",  x"d8", -- 1E80
         x"cd",  x"8d",  x"ce",  x"55",  x"cf",  x"95",  x"cd",  x"6d", -- 1E88
         x"cf",  x"64",  x"cd",  x"64",  x"cd",  x"23",  x"cd",  x"73", -- 1E90
         x"cd",  x"2c",  x"c9",  x"1f",  x"00",  x"96",  x"cb",  x"55", -- 1E98
         x"cf",  x"64",  x"cd",  x"98",  x"cc",  x"2c",  x"c9",  x"24", -- 1EA0
         x"00",  x"7c",  x"d0",  x"68",  x"c9",  x"0e",  x"00",  x"fa", -- 1EA8
         x"ca",  x"56",  x"ce",  x"55",  x"cf",  x"95",  x"cd",  x"50", -- 1EB0
         x"c9",  x"06",  x"00",  x"9a",  x"d0",  x"9a",  x"d0",  x"23", -- 1EB8
         x"cd",  x"81",  x"d6",  x"29",  x"d1",  x"f5",  x"d0",  x"64", -- 1EC0
         x"cd",  x"23",  x"cd",  x"74",  x"cc",  x"e5",  x"ca",  x"a8", -- 1EC8
         x"cb",  x"68",  x"c9",  x"c2",  x"ff",  x"09",  x"cd",  x"18", -- 1ED0
         x"cc",  x"84",  x"4c",  x"49",  x"53",  x"d4",  x"7f",  x"de", -- 1ED8
         x"d8",  x"cd",  x"47",  x"d2",  x"fa",  x"ca",  x"23",  x"cd", -- 1EE0
         x"5f",  x"cf",  x"95",  x"cd",  x"34",  x"d3",  x"06",  x"53", -- 1EE8
         x"43",  x"52",  x"20",  x"23",  x"20",  x"5e",  x"de",  x"8d", -- 1EF0
         x"ce",  x"99",  x"ce",  x"02",  x"da",  x"81",  x"ce",  x"21", -- 1EF8
         x"da",  x"56",  x"ce",  x"cb",  x"c9",  x"fa",  x"ca",  x"e7", -- 1F00
         x"c9",  x"2c",  x"c9",  x"03",  x"00",  x"3f",  x"de",  x"9a", -- 1F08
         x"d0",  x"e7",  x"c9",  x"5f",  x"cf",  x"64",  x"cd",  x"b3", -- 1F10
         x"da",  x"e5",  x"ca",  x"68",  x"c9",  x"0a",  x"00",  x"56", -- 1F18
         x"ce",  x"c3",  x"cf",  x"95",  x"cd",  x"2f",  x"cc",  x"7d", -- 1F20
         x"c9",  x"dc",  x"ff",  x"fa",  x"ca",  x"18",  x"cc",  x"85", -- 1F28
         x"49",  x"4e",  x"44",  x"45",  x"d8",  x"d9",  x"de",  x"d8", -- 1F30
         x"cd",  x"2c",  x"c9",  x"0c",  x"00",  x"a5",  x"ca",  x"fa", -- 1F38
         x"ca",  x"d6",  x"cf",  x"16",  x"cd",  x"cb",  x"c9",  x"fa", -- 1F40
         x"ca",  x"e7",  x"c9",  x"2c",  x"c9",  x"03",  x"00",  x"3f", -- 1F48
         x"de",  x"9a",  x"d0",  x"56",  x"ce",  x"e7",  x"c9",  x"b3", -- 1F50
         x"da",  x"e5",  x"ca",  x"68",  x"c9",  x"04",  x"00",  x"2f", -- 1F58
         x"cc",  x"7d",  x"c9",  x"e4",  x"ff",  x"18",  x"cc",  x"85", -- 1F60
         x"54",  x"52",  x"49",  x"41",  x"c4",  x"2f",  x"df",  x"d8", -- 1F68
         x"cd",  x"2c",  x"c9",  x"0c",  x"00",  x"a5",  x"ca",  x"2c", -- 1F70
         x"c9",  x"03",  x"00",  x"21",  x"da",  x"2c",  x"c9",  x"03", -- 1F78
         x"00",  x"02",  x"da",  x"2c",  x"c9",  x"03",  x"00",  x"fa", -- 1F80
         x"cc",  x"98",  x"cc",  x"16",  x"cd",  x"cb",  x"c9",  x"e7", -- 1F88
         x"c9",  x"a9",  x"d0",  x"68",  x"c9",  x"12",  x"00",  x"fa", -- 1F90
         x"ca",  x"e0",  x"de",  x"c3",  x"cf",  x"64",  x"cd",  x"74", -- 1F98
         x"cc",  x"68",  x"c9",  x"04",  x"00",  x"2f",  x"cc",  x"7d", -- 1FA0
         x"c9",  x"e6",  x"ff",  x"fa",  x"ca",  x"2c",  x"c9",  x"0f", -- 1FA8
         x"00",  x"c7",  x"da",  x"fa",  x"ca",  x"18",  x"cc",  x"85", -- 1FB0
         x"42",  x"55",  x"53",  x"49",  x"ce",  x"67",  x"df",  x"c1", -- 1FB8
         x"df",  x"d9",  x"e1",  x"4d",  x"ed",  x"78",  x"d9",  x"6f", -- 1FC0
         x"26",  x"00",  x"c3",  x"1a",  x"c9",  x"86",  x"42",  x"55", -- 1FC8
         x"53",  x"4f",  x"55",  x"d4",  x"b7",  x"df",  x"d8",  x"df", -- 1FD0
         x"d9",  x"e1",  x"d1",  x"4d",  x"ed",  x"59",  x"d9",  x"c3", -- 1FD8
         x"1b",  x"c9",  x"12",  x"00",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FF0
         x"cf",  x"57",  x"53",  x"d8",  x"bb",  x"a7",  x"64",  x"9e"  -- 1FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
