library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity caos_e is
    generic(
        ADDR_WIDTH   : integer := 13
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end caos_e;

architecture rtl of caos_e is
    type rom8192x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom8192x8 := (
         x"c3",  x"f6",  x"f0",  x"c3",  x"4f",  x"e6",  x"c3",  x"63", -- 0000
         x"e6",  x"c3",  x"db",  x"e6",  x"08",  x"fd",  x"c3",  x"a7", -- 0008
         x"f8",  x"7f",  x"7f",  x"42",  x"41",  x"53",  x"49",  x"43", -- 0010
         x"00",  x"cd",  x"2f",  x"e0",  x"c3",  x"0d",  x"c0",  x"7f", -- 0018
         x"7f",  x"52",  x"45",  x"42",  x"41",  x"53",  x"49",  x"43", -- 0020
         x"00",  x"cd",  x"2f",  x"e0",  x"c3",  x"8c",  x"c0",  x"db", -- 0028
         x"88",  x"f6",  x"80",  x"d3",  x"88",  x"dd",  x"7e",  x"04", -- 0030
         x"f6",  x"60",  x"d3",  x"86",  x"dd",  x"77",  x"04",  x"c9", -- 0038
         x"ed",  x"5b",  x"a0",  x"b7",  x"2a",  x"9c",  x"b7",  x"19", -- 0040
         x"cb",  x"24",  x"cb",  x"24",  x"cb",  x"24",  x"f5",  x"7d", -- 0048
         x"6c",  x"fe",  x"28",  x"30",  x"06",  x"f6",  x"80",  x"67", -- 0050
         x"f1",  x"a7",  x"c9",  x"f1",  x"37",  x"c9",  x"3a",  x"9e", -- 0058
         x"b7",  x"3d",  x"93",  x"d8",  x"3a",  x"9f",  x"b7",  x"3d", -- 0060
         x"92",  x"c9",  x"f5",  x"cd",  x"5e",  x"e0",  x"38",  x"eb", -- 0068
         x"3a",  x"9c",  x"b7",  x"83",  x"d5",  x"5f",  x"3a",  x"9d", -- 0070
         x"b7",  x"82",  x"87",  x"87",  x"87",  x"6f",  x"26",  x"00", -- 0078
         x"54",  x"29",  x"29",  x"19",  x"ed",  x"5b",  x"cb",  x"b7", -- 0080
         x"5f",  x"19",  x"d1",  x"f1",  x"a7",  x"c9",  x"f5",  x"e6", -- 0088
         x"c0",  x"4f",  x"f1",  x"f5",  x"e6",  x"07",  x"07",  x"07", -- 0090
         x"07",  x"b1",  x"4f",  x"f1",  x"0f",  x"0f",  x"0f",  x"e6", -- 0098
         x"07",  x"b1",  x"c9",  x"e5",  x"d5",  x"c5",  x"f5",  x"2a", -- 00A0
         x"9c",  x"b7",  x"19",  x"eb",  x"21",  x"a6",  x"b7",  x"87", -- 00A8
         x"30",  x"02",  x"2e",  x"aa",  x"d6",  x"40",  x"38",  x"04", -- 00B0
         x"fe",  x"80",  x"38",  x"04",  x"c6",  x"40",  x"2c",  x"2c", -- 00B8
         x"4e",  x"2c",  x"46",  x"87",  x"6f",  x"26",  x"00",  x"29", -- 00C0
         x"09",  x"7b",  x"fe",  x"28",  x"30",  x"56",  x"f6",  x"80", -- 00C8
         x"42",  x"57",  x"78",  x"87",  x"87",  x"87",  x"5f",  x"3a", -- 00D0
         x"a2",  x"b7",  x"cb",  x"57",  x"28",  x"0f",  x"4f",  x"06", -- 00D8
         x"08",  x"d5",  x"7e",  x"2f",  x"12",  x"23",  x"13",  x"10", -- 00E0
         x"f9",  x"79",  x"0f",  x"18",  x"14",  x"0f",  x"38",  x"12", -- 00E8
         x"d5",  x"ed",  x"a0",  x"ed",  x"a0",  x"ed",  x"a0",  x"ed", -- 00F0
         x"a0",  x"ed",  x"a0",  x"ed",  x"a0",  x"ed",  x"a0",  x"ed", -- 00F8
         x"a0",  x"d1",  x"0f",  x"38",  x"1f",  x"dd",  x"7e",  x"01", -- 0100
         x"67",  x"ee",  x"02",  x"f3",  x"d3",  x"84",  x"3a",  x"a3", -- 0108
         x"b7",  x"12",  x"13",  x"12",  x"13",  x"12",  x"13",  x"12", -- 0110
         x"13",  x"12",  x"13",  x"12",  x"13",  x"12",  x"13",  x"12", -- 0118
         x"7c",  x"d3",  x"84",  x"fb",  x"f1",  x"c1",  x"d1",  x"e1", -- 0120
         x"c9",  x"e5",  x"d5",  x"c5",  x"f5",  x"08",  x"f5",  x"79", -- 0128
         x"08",  x"3a",  x"9e",  x"b7",  x"e5",  x"d5",  x"ed",  x"a0", -- 0130
         x"ed",  x"a0",  x"ed",  x"a0",  x"ed",  x"a0",  x"ed",  x"a0", -- 0138
         x"ed",  x"a0",  x"ed",  x"a0",  x"ed",  x"a0",  x"ea",  x"36", -- 0140
         x"e1",  x"d1",  x"e1",  x"24",  x"14",  x"08",  x"4f",  x"08", -- 0148
         x"3d",  x"20",  x"e1",  x"08",  x"f1",  x"08",  x"18",  x"cc", -- 0150
         x"ed",  x"5b",  x"a0",  x"b7",  x"21",  x"a2",  x"b7",  x"cb", -- 0158
         x"66",  x"28",  x"22",  x"cb",  x"a6",  x"fe",  x"30",  x"d8", -- 0160
         x"fe",  x"3a",  x"30",  x"04",  x"d6",  x"30",  x"18",  x"0a", -- 0168
         x"fe",  x"41",  x"d8",  x"cb",  x"af",  x"fe",  x"5b",  x"d0", -- 0170
         x"d6",  x"37",  x"21",  x"df",  x"b7",  x"be",  x"d0",  x"87", -- 0178
         x"2a",  x"dd",  x"b7",  x"18",  x"0c",  x"fe",  x"20",  x"30", -- 0180
         x"19",  x"cb",  x"5e",  x"20",  x"15",  x"87",  x"2a",  x"b2", -- 0188
         x"b7",  x"4f",  x"06",  x"00",  x"09",  x"7e",  x"23",  x"66", -- 0190
         x"6f",  x"e9",  x"7b",  x"e6",  x"f8",  x"c6",  x"08",  x"5f", -- 0198
         x"18",  x"09",  x"cd",  x"6a",  x"e0",  x"d8",  x"77",  x"cd", -- 01A0
         x"a3",  x"e0",  x"1c",  x"3a",  x"9e",  x"b7",  x"3d",  x"bb", -- 01A8
         x"d0",  x"1e",  x"00",  x"14",  x"3a",  x"9f",  x"b7",  x"ba", -- 01B0
         x"c0",  x"2a",  x"a4",  x"b7",  x"e9",  x"2a",  x"99",  x"b7", -- 01B8
         x"e9",  x"7b",  x"a7",  x"28",  x"02",  x"1d",  x"c9",  x"7a", -- 01C0
         x"a7",  x"c8",  x"15",  x"3a",  x"9e",  x"b7",  x"3d",  x"5f", -- 01C8
         x"c9",  x"7a",  x"a7",  x"c8",  x"15",  x"c9",  x"21",  x"45", -- 01D0
         x"e2",  x"22",  x"a4",  x"b7",  x"c9",  x"21",  x"60",  x"e2", -- 01D8
         x"18",  x"f7",  x"cd",  x"c1",  x"e1",  x"d5",  x"cd",  x"6a", -- 01E0
         x"e0",  x"7e",  x"a7",  x"28",  x"29",  x"e5",  x"d5",  x"1c", -- 01E8
         x"cd",  x"6a",  x"e0",  x"30",  x"08",  x"1e",  x"00",  x"14", -- 01F0
         x"cd",  x"6a",  x"e0",  x"38",  x"10",  x"7e",  x"a7",  x"28", -- 01F8
         x"0c",  x"42",  x"4b",  x"d1",  x"e3",  x"77",  x"cd",  x"a3", -- 0200
         x"e0",  x"50",  x"59",  x"18",  x"e1",  x"d1",  x"e1",  x"36", -- 0208
         x"00",  x"3e",  x"20",  x"cd",  x"a3",  x"e0",  x"d1",  x"c9", -- 0210
         x"d5",  x"3e",  x"20",  x"cd",  x"6a",  x"e0",  x"46",  x"77", -- 0218
         x"cd",  x"a3",  x"e0",  x"78",  x"a7",  x"28",  x"0e",  x"1c", -- 0220
         x"cd",  x"6a",  x"e0",  x"30",  x"f1",  x"1e",  x"00",  x"14", -- 0228
         x"cd",  x"6a",  x"e0",  x"30",  x"e9",  x"d1",  x"c9",  x"3a", -- 0230
         x"9f",  x"b7",  x"16",  x"00",  x"f5",  x"cd",  x"aa",  x"e2", -- 0238
         x"f1",  x"14",  x"3d",  x"20",  x"f7",  x"16",  x"00",  x"1e", -- 0240
         x"00",  x"c9",  x"41",  x"55",  x"77",  x"2c",  x"77",  x"2c", -- 0248
         x"77",  x"2c",  x"77",  x"2c",  x"77",  x"2c",  x"77",  x"2c", -- 0250
         x"77",  x"2c",  x"77",  x"6a",  x"24",  x"10",  x"ec",  x"c9", -- 0258
         x"3a",  x"9e",  x"b7",  x"4f",  x"06",  x"00",  x"3a",  x"9f", -- 0260
         x"b7",  x"3d",  x"28",  x"3d",  x"d5",  x"f5",  x"11",  x"00", -- 0268
         x"00",  x"cd",  x"6a",  x"e0",  x"eb",  x"21",  x"28",  x"00", -- 0270
         x"19",  x"e5",  x"c5",  x"ed",  x"b0",  x"c1",  x"d1",  x"3d", -- 0278
         x"20",  x"f3",  x"f1",  x"87",  x"87",  x"87",  x"4f",  x"11", -- 0280
         x"00",  x"00",  x"42",  x"cd",  x"44",  x"e0",  x"eb",  x"2e", -- 0288
         x"08",  x"19",  x"3a",  x"a2",  x"b7",  x"1f",  x"1f",  x"38", -- 0290
         x"0b",  x"f5",  x"cd",  x"de",  x"e2",  x"cd",  x"29",  x"e1", -- 0298
         x"cd",  x"de",  x"e2",  x"f1",  x"17",  x"d4",  x"29",  x"e1", -- 02A0
         x"d1",  x"15",  x"1e",  x"00",  x"cd",  x"6a",  x"e0",  x"d8", -- 02A8
         x"3a",  x"9e",  x"b7",  x"47",  x"4f",  x"af",  x"77",  x"23", -- 02B0
         x"10",  x"fc",  x"cd",  x"44",  x"e0",  x"d8",  x"d5",  x"3a", -- 02B8
         x"a2",  x"b7",  x"0f",  x"5f",  x"38",  x"06",  x"af",  x"e5", -- 02C0
         x"cd",  x"4a",  x"e2",  x"e1",  x"cb",  x"0b",  x"38",  x"0c", -- 02C8
         x"cd",  x"de",  x"e2",  x"3a",  x"a3",  x"b7",  x"cd",  x"4a", -- 02D0
         x"e2",  x"cd",  x"de",  x"e2",  x"d1",  x"c9",  x"dd",  x"7e", -- 02D8
         x"01",  x"ee",  x"02",  x"f3",  x"dd",  x"77",  x"01",  x"d3", -- 02E0
         x"84",  x"fb",  x"c9",  x"01",  x"0f",  x"0a",  x"21",  x"30", -- 02E8
         x"00",  x"d5",  x"5c",  x"cd",  x"2e",  x"f9",  x"3e",  x"1e", -- 02F0
         x"cd",  x"e0",  x"f1",  x"3e",  x"03",  x"d3",  x"8c",  x"3e", -- 02F8
         x"10",  x"d1",  x"c3",  x"e0",  x"f1",  x"21",  x"30",  x"00", -- 0300
         x"d5",  x"5c",  x"cd",  x"2e",  x"f9",  x"d1",  x"c9",  x"21", -- 0308
         x"a3",  x"b7",  x"7e",  x"cd",  x"8e",  x"e0",  x"77",  x"c9", -- 0310
         x"7e",  x"c9",  x"dd",  x"7e",  x"08",  x"ee",  x"20",  x"dd", -- 0318
         x"77",  x"08",  x"c9",  x"21",  x"a2",  x"b7",  x"cb",  x"e6", -- 0320
         x"c9",  x"e5",  x"d5",  x"c5",  x"f5",  x"cd",  x"58",  x"e1", -- 0328
         x"ed",  x"53",  x"a0",  x"b7",  x"f1",  x"c1",  x"d1",  x"e1", -- 0330
         x"c9",  x"fb",  x"f5",  x"3e",  x"23",  x"d3",  x"8f",  x"dd", -- 0338
         x"36",  x"0d",  x"00",  x"18",  x"5e",  x"f5",  x"db",  x"8f", -- 0340
         x"f5",  x"3e",  x"a7",  x"d3",  x"8f",  x"3e",  x"8f",  x"d3", -- 0348
         x"8f",  x"f1",  x"fb",  x"b7",  x"28",  x"4d",  x"fe",  x"14", -- 0350
         x"38",  x"49",  x"fe",  x"78",  x"30",  x"45",  x"fe",  x"65", -- 0358
         x"30",  x"3d",  x"c6",  x"be",  x"38",  x"39",  x"e5",  x"d5", -- 0360
         x"dd",  x"7e",  x"0c",  x"1f",  x"ee",  x"01",  x"dd",  x"6e", -- 0368
         x"0e",  x"dd",  x"66",  x"0f",  x"16",  x"00",  x"5f",  x"19", -- 0370
         x"7e",  x"d1",  x"e1",  x"dd",  x"cb",  x"08",  x"7e",  x"20", -- 0378
         x"0a",  x"fe",  x"40",  x"38",  x"06",  x"fe",  x"80",  x"30", -- 0380
         x"02",  x"ee",  x"20",  x"dd",  x"be",  x"0d",  x"20",  x"1d", -- 0388
         x"f5",  x"3a",  x"e0",  x"b7",  x"dd",  x"be",  x"0a",  x"38", -- 0390
         x"11",  x"f1",  x"dd",  x"34",  x"0a",  x"18",  x"04",  x"dd", -- 0398
         x"cb",  x"0c",  x"1e",  x"db",  x"89",  x"d3",  x"89",  x"f1", -- 03A0
         x"ed",  x"4d",  x"f1",  x"18",  x"08",  x"dd",  x"36",  x"0a", -- 03A8
         x"00",  x"fe",  x"16",  x"28",  x"09",  x"dd",  x"77",  x"0d", -- 03B0
         x"dd",  x"cb",  x"08",  x"c6",  x"18",  x"e5",  x"dd",  x"7e", -- 03B8
         x"08",  x"ee",  x"80",  x"dd",  x"77",  x"08",  x"3e",  x"16", -- 03C0
         x"18",  x"eb",  x"b7",  x"dd",  x"cb",  x"08",  x"46",  x"c8", -- 03C8
         x"dd",  x"7e",  x"0d",  x"37",  x"c9",  x"cd",  x"ca",  x"e3", -- 03D0
         x"d0",  x"dd",  x"cb",  x"08",  x"86",  x"c9",  x"cd",  x"ca", -- 03D8
         x"e3",  x"d0",  x"fe",  x"03",  x"37",  x"c8",  x"a7",  x"c9", -- 03E0
         x"7f",  x"7f",  x"53",  x"57",  x"49",  x"54",  x"43",  x"48", -- 03E8
         x"01",  x"53",  x"cd",  x"04",  x"e4",  x"7d",  x"cd",  x"59", -- 03F0
         x"f3",  x"7c",  x"cd",  x"59",  x"f3",  x"7a",  x"cd",  x"76", -- 03F8
         x"f3",  x"c3",  x"6b",  x"f3",  x"26",  x"b8",  x"0e",  x"80", -- 0400
         x"45",  x"fe",  x"02",  x"30",  x"04",  x"56",  x"ed",  x"60", -- 0408
         x"c9",  x"72",  x"7d",  x"fe",  x"05",  x"38",  x"14",  x"ed", -- 0410
         x"51",  x"18",  x"f3",  x"e6",  x"f5",  x"cb",  x"42",  x"28", -- 0418
         x"5c",  x"cb",  x"cf",  x"cb",  x"4a",  x"28",  x"56",  x"cb", -- 0420
         x"df",  x"18",  x"52",  x"fe",  x"04",  x"38",  x"18",  x"dd", -- 0428
         x"7e",  x"04",  x"e6",  x"fc",  x"cb",  x"42",  x"28",  x"08", -- 0430
         x"cb",  x"c7",  x"cb",  x"4a",  x"28",  x"02",  x"cb",  x"cf", -- 0438
         x"dd",  x"77",  x"04",  x"d3",  x"86",  x"18",  x"38",  x"fe", -- 0440
         x"03",  x"38",  x"24",  x"db",  x"89",  x"e6",  x"9f",  x"cb", -- 0448
         x"42",  x"28",  x"08",  x"cb",  x"ef",  x"cb",  x"4a",  x"28", -- 0450
         x"02",  x"cb",  x"f7",  x"d3",  x"89",  x"dd",  x"7e",  x"01", -- 0458
         x"f6",  x"10",  x"cb",  x"52",  x"20",  x"02",  x"ee",  x"10", -- 0460
         x"d3",  x"84",  x"dd",  x"77",  x"01",  x"18",  x"10",  x"fe", -- 0468
         x"02",  x"38",  x"0f",  x"db",  x"88",  x"cb",  x"42",  x"cb", -- 0470
         x"bf",  x"28",  x"02",  x"cb",  x"ff",  x"d3",  x"88",  x"26", -- 0478
         x"ff",  x"c9",  x"fe",  x"01",  x"db",  x"88",  x"da",  x"1b", -- 0480
         x"e4",  x"cb",  x"42",  x"cb",  x"97",  x"28",  x"ee",  x"cb", -- 0488
         x"d7",  x"18",  x"ea",  x"7f",  x"7f",  x"4a",  x"55",  x"4d", -- 0490
         x"50",  x"01",  x"7d",  x"47",  x"0e",  x"80",  x"ed",  x"78", -- 0498
         x"3c",  x"ca",  x"61",  x"f3",  x"3e",  x"ff",  x"26",  x"b8", -- 04A0
         x"68",  x"77",  x"f3",  x"ed",  x"79",  x"db",  x"88",  x"e6", -- 04A8
         x"7e",  x"c3",  x"b4",  x"b7",  x"f3",  x"db",  x"88",  x"f6", -- 04B0
         x"40",  x"e6",  x"df",  x"d3",  x"88",  x"fb",  x"2a",  x"a4", -- 04B8
         x"b7",  x"22",  x"cf",  x"b7",  x"cd",  x"fd",  x"f1",  x"22", -- 04C0
         x"cd",  x"b7",  x"cd",  x"d6",  x"e1",  x"3e",  x"03",  x"d3", -- 04C8
         x"8c",  x"d3",  x"8d",  x"dd",  x"cb",  x"08",  x"8e",  x"18", -- 04D0
         x"28",  x"dd",  x"36",  x"02",  x"fe",  x"cd",  x"2b",  x"e5", -- 04D8
         x"2a",  x"cd",  x"b7",  x"22",  x"b9",  x"b7",  x"2a",  x"cf", -- 04E0
         x"b7",  x"22",  x"a4",  x"b7",  x"21",  x"80",  x"b7",  x"af", -- 04E8
         x"2d",  x"77",  x"20",  x"fc",  x"db",  x"88",  x"e6",  x"9f", -- 04F0
         x"d3",  x"88",  x"cd",  x"6b",  x"f3",  x"dd",  x"cb",  x"08", -- 04F8
         x"86",  x"dd",  x"cb",  x"01",  x"5e",  x"28",  x"06",  x"db", -- 0500
         x"89",  x"cb",  x"ff",  x"d3",  x"89",  x"dd",  x"cb",  x"08", -- 0508
         x"4e",  x"20",  x"fa",  x"3e",  x"47",  x"d3",  x"8e",  x"3e", -- 0510
         x"0c",  x"d3",  x"8e",  x"c9",  x"f3",  x"db",  x"88",  x"f6", -- 0518
         x"60",  x"cd",  x"bb",  x"e4",  x"dd",  x"36",  x"02",  x"00", -- 0520
         x"01",  x"00",  x"10",  x"dd",  x"34",  x"02",  x"f3",  x"3e", -- 0528
         x"87",  x"d3",  x"8d",  x"3e",  x"2f",  x"d3",  x"8d",  x"fb", -- 0530
         x"57",  x"5f",  x"cd",  x"80",  x"e5",  x"ed",  x"a1",  x"ea", -- 0538
         x"3a",  x"e5",  x"cd",  x"7e",  x"e5",  x"dd",  x"7e",  x"02", -- 0540
         x"cd",  x"6b",  x"e5",  x"dd",  x"6e",  x"05",  x"dd",  x"66", -- 0548
         x"06",  x"06",  x"80",  x"7e",  x"cd",  x"6b",  x"e5",  x"79", -- 0550
         x"86",  x"4f",  x"23",  x"10",  x"f6",  x"cd",  x"6b",  x"e5", -- 0558
         x"7a",  x"cd",  x"83",  x"e5",  x"5d",  x"54",  x"3e",  x"03", -- 0560
         x"d3",  x"8d",  x"c9",  x"c5",  x"4f",  x"06",  x"08",  x"cb", -- 0568
         x"09",  x"1e",  x"17",  x"d4",  x"80",  x"e5",  x"1e",  x"2f", -- 0570
         x"dc",  x"80",  x"e5",  x"10",  x"f2",  x"c1",  x"1e",  x"5d", -- 0578
         x"cd",  x"83",  x"e5",  x"dd",  x"72",  x"00",  x"dd",  x"7e", -- 0580
         x"00",  x"a7",  x"20",  x"fa",  x"53",  x"c9",  x"cd",  x"b4", -- 0588
         x"e4",  x"3e",  x"83",  x"d3",  x"8a",  x"e5",  x"d5",  x"06", -- 0590
         x"16",  x"dd",  x"36",  x"0d",  x"00",  x"cd",  x"1a",  x"e6", -- 0598
         x"38",  x"f5",  x"fe",  x"ba",  x"cd",  x"ed",  x"e5",  x"38", -- 05A0
         x"ee",  x"10",  x"f2",  x"06",  x"02",  x"af",  x"4f",  x"dd", -- 05A8
         x"77",  x"00",  x"cd",  x"2d",  x"e6",  x"fe",  x"5d",  x"30", -- 05B0
         x"f2",  x"10",  x"f2",  x"cd",  x"39",  x"e6",  x"38",  x"25", -- 05B8
         x"dd",  x"77",  x"02",  x"06",  x"80",  x"dd",  x"6e",  x"05", -- 05C0
         x"dd",  x"66",  x"06",  x"cd",  x"39",  x"e6",  x"38",  x"15", -- 05C8
         x"77",  x"dd",  x"7e",  x"0d",  x"86",  x"dd",  x"77",  x"0d", -- 05D0
         x"23",  x"10",  x"f0",  x"cd",  x"39",  x"e6",  x"38",  x"05", -- 05D8
         x"dd",  x"96",  x"0d",  x"c6",  x"ff",  x"d1",  x"e1",  x"f3", -- 05E0
         x"3e",  x"03",  x"d3",  x"8a",  x"fb",  x"db",  x"88",  x"cb", -- 05E8
         x"ef",  x"30",  x"02",  x"cb",  x"af",  x"d3",  x"88",  x"c9", -- 05F0
         x"f5",  x"3e",  x"87",  x"d3",  x"8d",  x"dd",  x"7e",  x"00", -- 05F8
         x"d3",  x"8d",  x"dd",  x"36",  x"00",  x"00",  x"18",  x"0e", -- 0600
         x"f5",  x"db",  x"8e",  x"dd",  x"77",  x"00",  x"3e",  x"07", -- 0608
         x"d3",  x"8e",  x"3e",  x"a3",  x"d3",  x"8e",  x"f1",  x"fb", -- 0610
         x"ed",  x"4d",  x"dd",  x"36",  x"00",  x"00",  x"db",  x"88", -- 0618
         x"d3",  x"88",  x"dd",  x"7e",  x"00",  x"b7",  x"28",  x"f6", -- 0620
         x"4f",  x"dd",  x"36",  x"00",  x"00",  x"db",  x"88",  x"d3", -- 0628
         x"88",  x"dd",  x"7e",  x"00",  x"b7",  x"28",  x"f6",  x"81", -- 0630
         x"c9",  x"11",  x"00",  x"08",  x"cd",  x"1a",  x"e6",  x"38", -- 0638
         x"03",  x"fe",  x"ba",  x"d8",  x"3f",  x"cb",  x"1b",  x"15", -- 0640
         x"20",  x"f2",  x"cd",  x"1a",  x"e6",  x"7b",  x"c9",  x"78", -- 0648
         x"d6",  x"09",  x"38",  x"4f",  x"fe",  x"1b",  x"30",  x"4b", -- 0650
         x"07",  x"4f",  x"06",  x"00",  x"eb",  x"21",  x"ba",  x"fd", -- 0658
         x"c3",  x"b7",  x"c8",  x"7e",  x"fe",  x"df",  x"d8",  x"fe", -- 0660
         x"e3",  x"d0",  x"fe",  x"e1",  x"ca",  x"97",  x"ea",  x"3a", -- 0668
         x"fd",  x"03",  x"a7",  x"20",  x"2e",  x"3c",  x"32",  x"fd", -- 0670
         x"03",  x"e5",  x"21",  x"a3",  x"b7",  x"cd",  x"95",  x"ec", -- 0678
         x"e1",  x"32",  x"7e",  x"03",  x"7e",  x"fe",  x"df",  x"28", -- 0680
         x"1d",  x"fe",  x"e2",  x"ca",  x"9b",  x"e6",  x"cd",  x"bd", -- 0688
         x"c8",  x"cd",  x"14",  x"eb",  x"7e",  x"fe",  x"3b",  x"28", -- 0690
         x"3d",  x"18",  x"08",  x"cd",  x"bd",  x"c8",  x"cd",  x"30", -- 0698
         x"eb",  x"18",  x"f1",  x"c3",  x"48",  x"c3",  x"cd",  x"bd", -- 06A0
         x"c8",  x"cd",  x"fa",  x"ea",  x"7e",  x"fe",  x"3b",  x"28", -- 06A8
         x"25",  x"cd",  x"cc",  x"c8",  x"2c",  x"fe",  x"e0",  x"20", -- 06B0
         x"ea",  x"cd",  x"bd",  x"c8",  x"cd",  x"14",  x"eb",  x"cd", -- 06B8
         x"cc",  x"c8",  x"3b",  x"cd",  x"03",  x"cb",  x"3a",  x"7e", -- 06C0
         x"03",  x"e5",  x"21",  x"a3",  x"b7",  x"cd",  x"91",  x"ec", -- 06C8
         x"e1",  x"c1",  x"c9",  x"c5",  x"18",  x"a3",  x"cd",  x"bd", -- 06D0
         x"c8",  x"18",  x"e8",  x"79",  x"fe",  x"62",  x"ca",  x"4b", -- 06D8
         x"ea",  x"fe",  x"6e",  x"ca",  x"c3",  x"ec",  x"fe",  x"7c", -- 06E0
         x"ca",  x"a1",  x"ed",  x"fe",  x"76",  x"ca",  x"c4",  x"ed", -- 06E8
         x"d6",  x"3e",  x"38",  x"af",  x"fe",  x"07",  x"30",  x"ab", -- 06F0
         x"eb",  x"01",  x"b2",  x"fd",  x"e1",  x"6f",  x"09",  x"4e", -- 06F8
         x"23",  x"66",  x"69",  x"e5",  x"eb",  x"c9",  x"cd",  x"cc", -- 0700
         x"c8",  x"28",  x"cd",  x"21",  x"d4",  x"f5",  x"cd",  x"d6", -- 0708
         x"c8",  x"cd",  x"3a",  x"cd",  x"cd",  x"db",  x"c8",  x"f1", -- 0710
         x"e5",  x"f5",  x"cd",  x"30",  x"d3",  x"23",  x"23",  x"5e", -- 0718
         x"23",  x"56",  x"c1",  x"c5",  x"f5",  x"d5",  x"4f",  x"af", -- 0720
         x"b9",  x"28",  x"0c",  x"b8",  x"28",  x"09",  x"79",  x"05", -- 0728
         x"28",  x"05",  x"81",  x"38",  x"2b",  x"10",  x"fb",  x"47", -- 0730
         x"0e",  x"00",  x"c5",  x"cd",  x"e1",  x"d1",  x"c1",  x"c1", -- 0738
         x"c5",  x"cd",  x"7e",  x"d1",  x"e1",  x"e3",  x"7c",  x"e1", -- 0740
         x"e3",  x"6f",  x"24",  x"25",  x"e5",  x"c5",  x"28",  x"07", -- 0748
         x"cd",  x"f2",  x"d2",  x"c1",  x"e1",  x"18",  x"f4",  x"c1", -- 0750
         x"e1",  x"d1",  x"cd",  x"02",  x"d3",  x"c3",  x"a9",  x"d1", -- 0758
         x"1e",  x"1c",  x"c3",  x"56",  x"c3",  x"e5",  x"21",  x"0a", -- 0760
         x"00",  x"22",  x"54",  x"03",  x"2a",  x"5f",  x"03",  x"f5", -- 0768
         x"e5",  x"23",  x"23",  x"7e",  x"23",  x"66",  x"6f",  x"22", -- 0770
         x"4e",  x"03",  x"22",  x"52",  x"03",  x"ed",  x"5b",  x"d7", -- 0778
         x"03",  x"1b",  x"1b",  x"e1",  x"e5",  x"7e",  x"23",  x"66", -- 0780
         x"6f",  x"cd",  x"89",  x"c6",  x"e3",  x"20",  x"f4",  x"d1", -- 0788
         x"23",  x"23",  x"7e",  x"23",  x"66",  x"6f",  x"22",  x"50", -- 0790
         x"03",  x"06",  x"04",  x"f1",  x"21",  x"4e",  x"03",  x"e3", -- 0798
         x"28",  x"20",  x"cd",  x"86",  x"c9",  x"f5",  x"7a",  x"b3", -- 07A0
         x"ca",  x"67",  x"c9",  x"f1",  x"e3",  x"73",  x"23",  x"72", -- 07A8
         x"23",  x"28",  x"0f",  x"f5",  x"05",  x"28",  x"07",  x"f1", -- 07B0
         x"e3",  x"cd",  x"d6",  x"c8",  x"18",  x"e2",  x"f1",  x"c2", -- 07B8
         x"69",  x"ea",  x"2a",  x"50",  x"03",  x"ed",  x"5b",  x"4e", -- 07C0
         x"03",  x"cd",  x"89",  x"c6",  x"da",  x"67",  x"c9",  x"2a", -- 07C8
         x"5f",  x"03",  x"cd",  x"be",  x"c4",  x"38",  x"04",  x"28", -- 07D0
         x"cf",  x"18",  x"f7",  x"e1",  x"c5",  x"ed",  x"5b",  x"50", -- 07D8
         x"03",  x"21",  x"00",  x"00",  x"22",  x"50",  x"03",  x"60", -- 07E0
         x"69",  x"4e",  x"23",  x"46",  x"78",  x"b1",  x"28",  x"b8", -- 07E8
         x"23",  x"7e",  x"23",  x"66",  x"6f",  x"cd",  x"89",  x"c6", -- 07F0
         x"2a",  x"50",  x"03",  x"23",  x"22",  x"50",  x"03",  x"20", -- 07F8
         x"e6",  x"23",  x"23",  x"29",  x"23",  x"ed",  x"5b",  x"d7", -- 0800
         x"03",  x"19",  x"38",  x"c0",  x"cd",  x"27",  x"c3",  x"22", -- 0808
         x"d7",  x"03",  x"af",  x"2b",  x"77",  x"2b",  x"77",  x"1b", -- 0810
         x"1b",  x"eb",  x"73",  x"23",  x"72",  x"23",  x"3d",  x"77", -- 0818
         x"23",  x"77",  x"23",  x"eb",  x"2a",  x"52",  x"03",  x"22", -- 0820
         x"4e",  x"03",  x"e1",  x"4e",  x"23",  x"46",  x"23",  x"c5", -- 0828
         x"01",  x"4e",  x"03",  x"7e",  x"12",  x"0a",  x"77",  x"23", -- 0830
         x"13",  x"03",  x"7e",  x"12",  x"0a",  x"77",  x"13",  x"2a", -- 0838
         x"4e",  x"03",  x"ed",  x"4b",  x"54",  x"03",  x"09",  x"22", -- 0840
         x"4e",  x"03",  x"2a",  x"50",  x"03",  x"2b",  x"7c",  x"b5", -- 0848
         x"22",  x"50",  x"03",  x"20",  x"d5",  x"12",  x"e1",  x"2a", -- 0850
         x"5f",  x"03",  x"e5",  x"e1",  x"4e",  x"23",  x"46",  x"23", -- 0858
         x"c5",  x"7e",  x"23",  x"a6",  x"3c",  x"28",  x"26",  x"23", -- 0860
         x"7e",  x"b7",  x"28",  x"ef",  x"fe",  x"88",  x"28",  x"2a", -- 0868
         x"fe",  x"8c",  x"28",  x"26",  x"fe",  x"8b",  x"28",  x"08", -- 0870
         x"fe",  x"d4",  x"28",  x"04",  x"fe",  x"a9",  x"20",  x"e7", -- 0878
         x"cd",  x"87",  x"c9",  x"7b",  x"b2",  x"c4",  x"ae",  x"e8", -- 0880
         x"c4",  x"e0",  x"e8",  x"18",  x"db",  x"2b",  x"22",  x"d7", -- 0888
         x"03",  x"2b",  x"77",  x"2b",  x"77",  x"e1",  x"e1",  x"c3", -- 0890
         x"8a",  x"c4",  x"cd",  x"87",  x"c9",  x"7b",  x"b2",  x"28", -- 0898
         x"c7",  x"cd",  x"ae",  x"e8",  x"c4",  x"e0",  x"e8",  x"7e", -- 08A0
         x"fe",  x"2c",  x"20",  x"bc",  x"18",  x"ec",  x"e5",  x"d5", -- 08A8
         x"11",  x"ff",  x"ff",  x"cd",  x"bb",  x"c4",  x"d1",  x"03", -- 08B0
         x"03",  x"03",  x"03",  x"60",  x"69",  x"ed",  x"4b",  x"52", -- 08B8
         x"03",  x"7e",  x"23",  x"e5",  x"b6",  x"28",  x"16",  x"7e", -- 08C0
         x"2b",  x"6e",  x"67",  x"cd",  x"89",  x"c6",  x"28",  x"0a", -- 08C8
         x"2a",  x"54",  x"03",  x"09",  x"44",  x"4d",  x"e1",  x"23", -- 08D0
         x"18",  x"e7",  x"3e",  x"ff",  x"b7",  x"e1",  x"e1",  x"c9", -- 08D8
         x"c5",  x"eb",  x"2a",  x"d7",  x"03",  x"ed",  x"52",  x"e5", -- 08E0
         x"c1",  x"62",  x"6b",  x"1b",  x"1a",  x"fe",  x"2c",  x"28", -- 08E8
         x"0b",  x"fe",  x"3a",  x"30",  x"07",  x"c5",  x"d5",  x"ed", -- 08F0
         x"b0",  x"d1",  x"18",  x"ec",  x"eb",  x"d1",  x"e5",  x"c5", -- 08F8
         x"af",  x"06",  x"98",  x"cd",  x"ae",  x"d6",  x"cd",  x"34", -- 0900
         x"d8",  x"c1",  x"d1",  x"23",  x"13",  x"7e",  x"b7",  x"28", -- 0908
         x"0f",  x"c5",  x"e5",  x"eb",  x"09",  x"54",  x"5d",  x"2b", -- 0910
         x"ed",  x"b8",  x"e1",  x"ed",  x"a0",  x"c1",  x"18",  x"ed", -- 0918
         x"d5",  x"ed",  x"5b",  x"5f",  x"03",  x"cd",  x"93",  x"c4", -- 0920
         x"23",  x"7e",  x"23",  x"b6",  x"20",  x"fa",  x"eb",  x"73", -- 0928
         x"23",  x"72",  x"13",  x"13",  x"ed",  x"53",  x"d7",  x"03", -- 0930
         x"e1",  x"54",  x"5d",  x"7e",  x"b7",  x"23",  x"20",  x"fb", -- 0938
         x"c1",  x"e3",  x"c5",  x"eb",  x"c9",  x"c8",  x"cd",  x"86", -- 0940
         x"c9",  x"ca",  x"42",  x"c4",  x"cd",  x"d6",  x"c8",  x"d5", -- 0948
         x"cd",  x"86",  x"c9",  x"e1",  x"c0",  x"eb",  x"e5",  x"cd", -- 0950
         x"bb",  x"c4",  x"d2",  x"4d",  x"c4",  x"d1",  x"f5",  x"c5", -- 0958
         x"cd",  x"be",  x"c4",  x"d2",  x"4d",  x"c4",  x"c1",  x"c3", -- 0960
         x"50",  x"c4",  x"cd",  x"be",  x"c8",  x"20",  x"0f",  x"cd", -- 0968
         x"ca",  x"e3",  x"30",  x"fb",  x"fe",  x"03",  x"c8",  x"fe", -- 0970
         x"0a",  x"20",  x"f4",  x"c3",  x"e4",  x"dd",  x"cd",  x"21", -- 0978
         x"d4",  x"4f",  x"3e",  x"10",  x"1e",  x"14",  x"cd",  x"15", -- 0980
         x"f0",  x"c5",  x"cd",  x"ca",  x"e3",  x"c1",  x"30",  x"0a", -- 0988
         x"fe",  x"03",  x"c8",  x"fe",  x"0a",  x"20",  x"03",  x"c3", -- 0990
         x"e4",  x"dd",  x"0d",  x"20",  x"e5",  x"c9",  x"06",  x"01", -- 0998
         x"cd",  x"be",  x"c8",  x"28",  x"04",  x"cd",  x"21",  x"d4", -- 09A0
         x"47",  x"3e",  x"07",  x"1e",  x"00",  x"cd",  x"15",  x"f0", -- 09A8
         x"10",  x"f7",  x"c9",  x"cd",  x"be",  x"c8",  x"28",  x"65", -- 09B0
         x"e5",  x"cd",  x"21",  x"d4",  x"e3",  x"21",  x"f6",  x"b9", -- 09B8
         x"cd",  x"91",  x"ec",  x"23",  x"e3",  x"cd",  x"d6",  x"c8", -- 09C0
         x"cd",  x"21",  x"d4",  x"e3",  x"cd",  x"91",  x"ec",  x"23", -- 09C8
         x"e3",  x"cd",  x"d6",  x"c8",  x"cd",  x"21",  x"d4",  x"e3", -- 09D0
         x"cd",  x"91",  x"ec",  x"e3",  x"cd",  x"d6",  x"c8",  x"cd", -- 09D8
         x"21",  x"d4",  x"e3",  x"57",  x"cd",  x"18",  x"f0",  x"fe", -- 09E0
         x"28",  x"30",  x"4d",  x"3a",  x"f8",  x"b9",  x"5f",  x"fe", -- 09E8
         x"28",  x"30",  x"45",  x"7a",  x"93",  x"38",  x"41",  x"3c", -- 09F0
         x"32",  x"9e",  x"b7",  x"7b",  x"32",  x"9c",  x"b7",  x"3a", -- 09F8
         x"f7",  x"b9",  x"fe",  x"20",  x"30",  x"32",  x"57",  x"3a", -- 0A00
         x"f6",  x"b9",  x"fe",  x"20",  x"30",  x"2a",  x"5f",  x"7a", -- 0A08
         x"93",  x"38",  x"25",  x"3c",  x"32",  x"9f",  x"b7",  x"7b", -- 0A10
         x"32",  x"9d",  x"b7",  x"18",  x"10",  x"e5",  x"cd",  x"18", -- 0A18
         x"f0",  x"21",  x"00",  x"01",  x"22",  x"9c",  x"b7",  x"21", -- 0A20
         x"28",  x"1e",  x"22",  x"9e",  x"b7",  x"21",  x"00",  x"00", -- 0A28
         x"22",  x"a0",  x"b7",  x"cd",  x"1b",  x"f0",  x"e1",  x"c9", -- 0A30
         x"cd",  x"1b",  x"f0",  x"18",  x"2c",  x"e5",  x"21",  x"81", -- 0A38
         x"b7",  x"af",  x"cd",  x"91",  x"ec",  x"e1",  x"1e",  x"10", -- 0A40
         x"c3",  x"15",  x"f0",  x"cd",  x"e1",  x"cd",  x"e3",  x"11", -- 0A48
         x"f3",  x"cd",  x"d5",  x"cd",  x"6f",  x"c9",  x"e5",  x"21", -- 0A50
         x"00",  x"80",  x"19",  x"38",  x"03",  x"3e",  x"bf",  x"bc", -- 0A58
         x"38",  x"07",  x"cd",  x"95",  x"ec",  x"e1",  x"c3",  x"e9", -- 0A60
         x"d3",  x"c3",  x"48",  x"c3",  x"cd",  x"6c",  x"c9",  x"d5", -- 0A68
         x"cd",  x"d6",  x"c8",  x"cd",  x"21",  x"d4",  x"e3",  x"11", -- 0A70
         x"00",  x"80",  x"19",  x"38",  x"e3",  x"57",  x"3e",  x"bf", -- 0A78
         x"bc",  x"38",  x"dd",  x"7a",  x"cd",  x"91",  x"ec",  x"e1", -- 0A80
         x"c9",  x"cd",  x"21",  x"d4",  x"0f",  x"0f",  x"0f",  x"e6", -- 0A88
         x"60",  x"4f",  x"06",  x"9f",  x"c3",  x"53",  x"f9",  x"3a", -- 0A90
         x"fd",  x"03",  x"cb",  x"4f",  x"cb",  x"cf",  x"32",  x"fd", -- 0A98
         x"03",  x"20",  x"c6",  x"d5",  x"e5",  x"cd",  x"18",  x"f0", -- 0AA0
         x"21",  x"9c",  x"b7",  x"22",  x"f6",  x"b9",  x"11",  x"ec", -- 0AA8
         x"b9",  x"01",  x"06",  x"00",  x"ed",  x"b0",  x"21",  x"00", -- 0AB0
         x"00",  x"22",  x"9c",  x"b7",  x"21",  x"28",  x"20",  x"22", -- 0AB8
         x"9e",  x"b7",  x"cd",  x"1b",  x"f0",  x"e1",  x"cd",  x"42", -- 0AC0
         x"eb",  x"cd",  x"db",  x"c8",  x"cd",  x"cc",  x"c8",  x"3b", -- 0AC8
         x"7e",  x"fe",  x"df",  x"38",  x"1d",  x"fe",  x"e3",  x"30", -- 0AD0
         x"19",  x"cd",  x"d3",  x"e6",  x"e5",  x"cd",  x"18",  x"f0", -- 0AD8
         x"21",  x"ec",  x"b9",  x"11",  x"9c",  x"b7",  x"01",  x"06", -- 0AE0
         x"00",  x"ed",  x"b0",  x"cd",  x"1b",  x"f0",  x"e1",  x"d1", -- 0AE8
         x"c1",  x"c9",  x"cd",  x"03",  x"cb",  x"18",  x"e5",  x"c3", -- 0AF0
         x"48",  x"c3",  x"cd",  x"21",  x"d4",  x"fe",  x"20",  x"30", -- 0AF8
         x"f6",  x"cb",  x"27",  x"cb",  x"27",  x"cb",  x"27",  x"57", -- 0B00
         x"e5",  x"21",  x"a3",  x"b7",  x"cd",  x"95",  x"ec",  x"e1", -- 0B08
         x"e6",  x"07",  x"18",  x"12",  x"cd",  x"21",  x"d4",  x"fe", -- 0B10
         x"08",  x"30",  x"dc",  x"57",  x"e5",  x"21",  x"a3",  x"b7", -- 0B18
         x"cd",  x"95",  x"ec",  x"e1",  x"e6",  x"f8",  x"b2",  x"e5", -- 0B20
         x"21",  x"a3",  x"b7",  x"cd",  x"91",  x"ec",  x"e1",  x"c9", -- 0B28
         x"cd",  x"be",  x"c8",  x"28",  x"c2",  x"cd",  x"fa",  x"ea", -- 0B30
         x"cd",  x"be",  x"c8",  x"c8",  x"cd",  x"d6",  x"c8",  x"18", -- 0B38
         x"d3",  x"c9",  x"cd",  x"bd",  x"c8",  x"cd",  x"cc",  x"c8", -- 0B40
         x"28",  x"cd",  x"21",  x"d4",  x"57",  x"e5",  x"21",  x"9f", -- 0B48
         x"b7",  x"cd",  x"95",  x"ec",  x"e1",  x"3d",  x"ba",  x"38", -- 0B50
         x"9e",  x"cd",  x"d6",  x"c8",  x"d5",  x"cd",  x"21",  x"d4", -- 0B58
         x"d1",  x"4f",  x"e5",  x"21",  x"9e",  x"b7",  x"cd",  x"95", -- 0B60
         x"ec",  x"e1",  x"3d",  x"b9",  x"38",  x"89",  x"79",  x"e5", -- 0B68
         x"21",  x"a0",  x"b7",  x"cd",  x"91",  x"ec",  x"7a",  x"23", -- 0B70
         x"cd",  x"91",  x"ec",  x"e1",  x"c9",  x"e5",  x"cd",  x"ca", -- 0B78
         x"e3",  x"30",  x"0f",  x"3e",  x"01",  x"cd",  x"7b",  x"d1", -- 0B80
         x"cd",  x"e4",  x"dd",  x"2a",  x"c2",  x"03",  x"77",  x"c3", -- 0B88
         x"a9",  x"d1",  x"af",  x"cd",  x"7b",  x"d1",  x"18",  x"f7", -- 0B90
         x"cd",  x"21",  x"d4",  x"e5",  x"21",  x"82",  x"b7",  x"06", -- 0B98
         x"04",  x"cd",  x"91",  x"ec",  x"23",  x"e3",  x"05",  x"28", -- 0BA0
         x"0b",  x"c5",  x"cd",  x"d6",  x"c8",  x"cd",  x"21",  x"d4", -- 0BA8
         x"c1",  x"e3",  x"18",  x"ed",  x"cd",  x"be",  x"c8",  x"28", -- 0BB0
         x"1c",  x"cd",  x"d6",  x"c8",  x"cd",  x"21",  x"d4",  x"e3", -- 0BB8
         x"cd",  x"91",  x"ec",  x"23",  x"e3",  x"cd",  x"be",  x"c8", -- 0BC0
         x"28",  x"0b",  x"cd",  x"d6",  x"c8",  x"cd",  x"21",  x"d4", -- 0BC8
         x"e3",  x"cd",  x"91",  x"ec",  x"e3",  x"1e",  x"35",  x"c1", -- 0BD0
         x"c3",  x"15",  x"f0",  x"06",  x"01",  x"c5",  x"cd",  x"6c", -- 0BD8
         x"c9",  x"e5",  x"7b",  x"21",  x"d3",  x"b7",  x"cd",  x"91", -- 0BE0
         x"ec",  x"7a",  x"23",  x"cd",  x"91",  x"ec",  x"e3",  x"cd", -- 0BE8
         x"d6",  x"c8",  x"cd",  x"21",  x"d4",  x"e3",  x"23",  x"cd", -- 0BF0
         x"91",  x"ec",  x"e1",  x"cd",  x"10",  x"ec",  x"1e",  x"30", -- 0BF8
         x"c1",  x"05",  x"28",  x"01",  x"1d",  x"cd",  x"15",  x"f0", -- 0C00
         x"da",  x"69",  x"ea",  x"c9",  x"06",  x"00",  x"18",  x"cd", -- 0C08
         x"cd",  x"be",  x"c8",  x"c8",  x"cd",  x"d6",  x"c8",  x"cd", -- 0C10
         x"21",  x"d4",  x"e5",  x"21",  x"d6",  x"b7",  x"17",  x"17", -- 0C18
         x"17",  x"c3",  x"78",  x"eb",  x"cd",  x"36",  x"cd",  x"cd", -- 0C20
         x"d6",  x"c8",  x"e5",  x"cd",  x"30",  x"d3",  x"28",  x"38", -- 0C28
         x"47",  x"23",  x"23",  x"5e",  x"23",  x"56",  x"e1",  x"d5", -- 0C30
         x"c5",  x"cd",  x"3a",  x"cd",  x"cd",  x"db",  x"c8",  x"c1", -- 0C38
         x"d1",  x"e5",  x"d5",  x"c5",  x"cd",  x"30",  x"d3",  x"28", -- 0C40
         x"1f",  x"23",  x"23",  x"4e",  x"23",  x"66",  x"69",  x"c1", -- 0C48
         x"4f",  x"d1",  x"e5",  x"c5",  x"d5",  x"1a",  x"be",  x"28", -- 0C50
         x"12",  x"23",  x"0d",  x"20",  x"f9",  x"af",  x"e1",  x"e1", -- 0C58
         x"e1",  x"11",  x"f3",  x"cd",  x"d5",  x"c3",  x"c0",  x"d0", -- 0C60
         x"c3",  x"67",  x"c9",  x"23",  x"e5",  x"2b",  x"23",  x"0d", -- 0C68
         x"28",  x"0e",  x"13",  x"05",  x"28",  x"11",  x"1a",  x"be", -- 0C70
         x"28",  x"f4",  x"e1",  x"d1",  x"c1",  x"0d",  x"18",  x"d3", -- 0C78
         x"13",  x"05",  x"e1",  x"20",  x"d8",  x"18",  x"01",  x"e1", -- 0C80
         x"d1",  x"d1",  x"d1",  x"a7",  x"ed",  x"52",  x"7d",  x"18", -- 0C88
         x"d0",  x"1e",  x"28",  x"18",  x"10",  x"1e",  x"29",  x"18", -- 0C90
         x"0c",  x"cd",  x"21",  x"d4",  x"a7",  x"28",  x"56",  x"fe", -- 0C98
         x"0d",  x"30",  x"52",  x"1e",  x"39",  x"c3",  x"15",  x"f0", -- 0CA0
         x"1e",  x"3a",  x"18",  x"f9",  x"cd",  x"21",  x"d4",  x"f5", -- 0CA8
         x"cd",  x"d6",  x"c8",  x"cd",  x"21",  x"d4",  x"57",  x"f1", -- 0CB0
         x"e5",  x"6f",  x"3e",  x"02",  x"1e",  x"26",  x"cd",  x"15", -- 0CB8
         x"f0",  x"e1",  x"c9",  x"cd",  x"e1",  x"cd",  x"e3",  x"11", -- 0CC0
         x"f3",  x"cd",  x"d5",  x"cd",  x"6f",  x"c9",  x"e5",  x"7b", -- 0CC8
         x"21",  x"d3",  x"b7",  x"cd",  x"91",  x"ec",  x"7a",  x"23", -- 0CD0
         x"cd",  x"91",  x"ec",  x"1e",  x"2f",  x"cd",  x"15",  x"f0", -- 0CD8
         x"06",  x"00",  x"28",  x"0c",  x"23",  x"23",  x"cd",  x"91", -- 0CE0
         x"ec",  x"1e",  x"30",  x"cd",  x"15",  x"f0",  x"06",  x"01", -- 0CE8
         x"78",  x"e1",  x"c3",  x"e9",  x"d3",  x"c3",  x"48",  x"c3", -- 0CF0
         x"0e",  x"00",  x"7e",  x"fe",  x"49",  x"28",  x"05",  x"0c", -- 0CF8
         x"fe",  x"4f",  x"20",  x"f1",  x"c5",  x"23",  x"7e",  x"fe", -- 0D00
         x"23",  x"20",  x"ea",  x"23",  x"cd",  x"21",  x"d4",  x"e6", -- 0D08
         x"03",  x"c1",  x"c8",  x"e5",  x"17",  x"81",  x"f5",  x"3d", -- 0D10
         x"06",  x"00",  x"37",  x"cb",  x"10",  x"3d",  x"20",  x"fb", -- 0D18
         x"21",  x"07",  x"03",  x"7e",  x"a8",  x"77",  x"f1",  x"e1", -- 0D20
         x"cb",  x"f7",  x"d5",  x"5f",  x"16",  x"03",  x"cd",  x"0e", -- 0D28
         x"e0",  x"d1",  x"c9",  x"ed",  x"5f",  x"32",  x"1d",  x"03", -- 0D30
         x"c9",  x"7e",  x"23",  x"fe",  x"49",  x"28",  x"19",  x"fe", -- 0D38
         x"4f",  x"20",  x"c6",  x"cd",  x"25",  x"de",  x"cd",  x"c8", -- 0D40
         x"dd",  x"c8",  x"3e",  x"d5",  x"cd",  x"b2",  x"dc",  x"21", -- 0D48
         x"ea",  x"03",  x"af",  x"cd",  x"d5",  x"dd",  x"e1",  x"c9", -- 0D50
         x"cd",  x"5f",  x"de",  x"3a",  x"09",  x"03",  x"e6",  x"03", -- 0D58
         x"c8",  x"3e",  x"d5",  x"cd",  x"b2",  x"dc",  x"21",  x"ea", -- 0D60
         x"03",  x"cd",  x"e4",  x"dd",  x"e1",  x"c9",  x"01",  x"3e", -- 0D68
         x"04",  x"18",  x"03",  x"01",  x"3f",  x"03",  x"c5",  x"cd", -- 0D70
         x"6c",  x"c9",  x"c1",  x"c5",  x"e5",  x"21",  x"82",  x"b7", -- 0D78
         x"7b",  x"cd",  x"91",  x"ec",  x"23",  x"7a",  x"cd",  x"91", -- 0D80
         x"ec",  x"23",  x"05",  x"28",  x"0c",  x"e3",  x"c5",  x"cd", -- 0D88
         x"d6",  x"c8",  x"cd",  x"6c",  x"c9",  x"c1",  x"e3",  x"18", -- 0D90
         x"e7",  x"e1",  x"cd",  x"10",  x"ec",  x"d1",  x"c3",  x"15", -- 0D98
         x"f0",  x"cd",  x"e1",  x"cd",  x"e3",  x"11",  x"f3",  x"cd", -- 0DA0
         x"d5",  x"cd",  x"24",  x"d4",  x"e5",  x"a7",  x"3e",  x"00", -- 0DA8
         x"20",  x"06",  x"21",  x"9d",  x"b7",  x"cd",  x"95",  x"ec", -- 0DB0
         x"47",  x"21",  x"a1",  x"b7",  x"cd",  x"95",  x"ec",  x"80", -- 0DB8
         x"e1",  x"c3",  x"e9",  x"d3",  x"e3",  x"3e",  x"01",  x"cd", -- 0DC0
         x"7b",  x"d1",  x"cd",  x"18",  x"f0",  x"ed",  x"5b",  x"a0", -- 0DC8
         x"b7",  x"cd",  x"6a",  x"e0",  x"7e",  x"cd",  x"1b",  x"f0", -- 0DD0
         x"c3",  x"8b",  x"eb",  x"9a",  x"e1",  x"6e",  x"f9",  x"7f", -- 0DD8
         x"f9",  x"8c",  x"f9",  x"9b",  x"f9",  x"8d",  x"f8",  x"9f", -- 0DE0
         x"f8",  x"aa",  x"f9",  x"0f",  x"e3",  x"b2",  x"f9",  x"b9", -- 0DE8
         x"f9",  x"00",  x"03",  x"c0",  x"20",  x"99",  x"c1",  x"00", -- 0DF0
         x"00",  x"4c",  x"58",  x"33",  x"00",  x"00",  x"00",  x"42", -- 0DF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0E00
         x"30",  x"30",  x"30",  x"30",  x"30",  x"00",  x"30",  x"00", -- 0E08
         x"77",  x"33",  x"66",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0E10
         x"36",  x"36",  x"fe",  x"6c",  x"fe",  x"d8",  x"d8",  x"00", -- 0E18
         x"18",  x"3e",  x"6c",  x"3e",  x"1b",  x"1b",  x"7e",  x"18", -- 0E20
         x"00",  x"c6",  x"cc",  x"18",  x"30",  x"66",  x"c6",  x"00", -- 0E28
         x"38",  x"6c",  x"38",  x"76",  x"dc",  x"cc",  x"76",  x"00", -- 0E30
         x"1c",  x"0c",  x"18",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0E38
         x"18",  x"30",  x"60",  x"60",  x"60",  x"30",  x"18",  x"00", -- 0E40
         x"60",  x"30",  x"18",  x"18",  x"18",  x"30",  x"60",  x"00", -- 0E48
         x"00",  x"66",  x"3c",  x"ff",  x"3c",  x"66",  x"00",  x"00", -- 0E50
         x"00",  x"30",  x"30",  x"fc",  x"30",  x"30",  x"00",  x"00", -- 0E58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"1c",  x"0c",  x"18", -- 0E60
         x"00",  x"00",  x"00",  x"fe",  x"00",  x"00",  x"00",  x"00", -- 0E68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"30",  x"30",  x"00", -- 0E70
         x"06",  x"0c",  x"18",  x"30",  x"60",  x"c0",  x"80",  x"00", -- 0E78
         x"7c",  x"c6",  x"ce",  x"de",  x"f6",  x"e6",  x"7c",  x"00", -- 0E80
         x"30",  x"70",  x"30",  x"30",  x"30",  x"30",  x"fc",  x"00", -- 0E88
         x"78",  x"cc",  x"0c",  x"38",  x"60",  x"cc",  x"fc",  x"00", -- 0E90
         x"fc",  x"18",  x"30",  x"78",  x"0c",  x"cc",  x"78",  x"00", -- 0E98
         x"1c",  x"3c",  x"6c",  x"cc",  x"fe",  x"0c",  x"1e",  x"00", -- 0EA0
         x"fc",  x"c0",  x"f8",  x"0c",  x"0c",  x"cc",  x"78",  x"00", -- 0EA8
         x"38",  x"60",  x"c0",  x"f8",  x"cc",  x"cc",  x"78",  x"00", -- 0EB0
         x"fc",  x"cc",  x"0c",  x"18",  x"30",  x"30",  x"30",  x"00", -- 0EB8
         x"78",  x"cc",  x"cc",  x"78",  x"cc",  x"cc",  x"78",  x"00", -- 0EC0
         x"78",  x"cc",  x"cc",  x"7c",  x"0c",  x"18",  x"70",  x"00", -- 0EC8
         x"00",  x"00",  x"30",  x"30",  x"00",  x"30",  x"30",  x"00", -- 0ED0
         x"00",  x"00",  x"30",  x"30",  x"00",  x"30",  x"30",  x"60", -- 0ED8
         x"18",  x"30",  x"60",  x"c0",  x"60",  x"30",  x"18",  x"00", -- 0EE0
         x"00",  x"00",  x"fc",  x"00",  x"fc",  x"00",  x"00",  x"00", -- 0EE8
         x"60",  x"30",  x"18",  x"0c",  x"18",  x"30",  x"60",  x"00", -- 0EF0
         x"78",  x"cc",  x"0c",  x"18",  x"30",  x"00",  x"30",  x"00", -- 0EF8
         x"7c",  x"c6",  x"de",  x"de",  x"de",  x"c0",  x"78",  x"00", -- 0F00
         x"30",  x"78",  x"cc",  x"cc",  x"fc",  x"cc",  x"cc",  x"00", -- 0F08
         x"fc",  x"66",  x"66",  x"7c",  x"66",  x"66",  x"fc",  x"00", -- 0F10
         x"3c",  x"66",  x"c0",  x"c0",  x"c0",  x"66",  x"3c",  x"00", -- 0F18
         x"f8",  x"6c",  x"66",  x"66",  x"66",  x"6c",  x"f8",  x"00", -- 0F20
         x"fe",  x"62",  x"68",  x"78",  x"68",  x"62",  x"fe",  x"00", -- 0F28
         x"fe",  x"62",  x"68",  x"78",  x"68",  x"60",  x"f0",  x"00", -- 0F30
         x"3c",  x"66",  x"c0",  x"c0",  x"ce",  x"66",  x"3c",  x"00", -- 0F38
         x"cc",  x"cc",  x"cc",  x"fc",  x"cc",  x"cc",  x"cc",  x"00", -- 0F40
         x"78",  x"30",  x"30",  x"30",  x"30",  x"30",  x"78",  x"00", -- 0F48
         x"1e",  x"0c",  x"0c",  x"0c",  x"cc",  x"cc",  x"78",  x"00", -- 0F50
         x"e6",  x"66",  x"6c",  x"70",  x"6c",  x"66",  x"e6",  x"00", -- 0F58
         x"f0",  x"60",  x"60",  x"60",  x"62",  x"66",  x"fe",  x"00", -- 0F60
         x"c6",  x"ee",  x"fe",  x"d6",  x"c6",  x"c6",  x"c6",  x"00", -- 0F68
         x"c6",  x"e6",  x"f6",  x"de",  x"ce",  x"c6",  x"c6",  x"00", -- 0F70
         x"38",  x"6c",  x"c6",  x"c6",  x"c6",  x"6c",  x"38",  x"00", -- 0F78
         x"fc",  x"66",  x"66",  x"7c",  x"60",  x"60",  x"f0",  x"00", -- 0F80
         x"78",  x"cc",  x"cc",  x"cc",  x"dc",  x"78",  x"1c",  x"00", -- 0F88
         x"fc",  x"66",  x"66",  x"7c",  x"6c",  x"66",  x"e6",  x"00", -- 0F90
         x"7c",  x"c6",  x"f0",  x"3c",  x"0e",  x"c6",  x"7c",  x"00", -- 0F98
         x"fc",  x"b4",  x"30",  x"30",  x"30",  x"30",  x"78",  x"00", -- 0FA0
         x"cc",  x"cc",  x"cc",  x"cc",  x"cc",  x"cc",  x"78",  x"00", -- 0FA8
         x"cc",  x"cc",  x"cc",  x"78",  x"78",  x"30",  x"30",  x"00", -- 0FB0
         x"c6",  x"c6",  x"c6",  x"d6",  x"fe",  x"ee",  x"c6",  x"00", -- 0FB8
         x"c6",  x"c6",  x"6c",  x"38",  x"6c",  x"c6",  x"c6",  x"00", -- 0FC0
         x"cc",  x"cc",  x"cc",  x"78",  x"30",  x"30",  x"78",  x"00", -- 0FC8
         x"fe",  x"c6",  x"8c",  x"18",  x"32",  x"66",  x"fe",  x"00", -- 0FD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FD8
         x"18",  x"18",  x"18",  x"18",  x"18",  x"18",  x"18",  x"00", -- 0FE0
         x"00",  x"fe",  x"06",  x"06",  x"00",  x"00",  x"00",  x"00", -- 0FE8
         x"10",  x"38",  x"6c",  x"c6",  x"00",  x"00",  x"00",  x"00", -- 0FF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"ff", -- 0FF8
         x"c3",  x"bf",  x"f0",  x"c3",  x"47",  x"f0",  x"c3",  x"63", -- 1000
         x"f0",  x"c3",  x"77",  x"f0",  x"c3",  x"33",  x"f0",  x"c3", -- 1008
         x"b0",  x"f0",  x"c3",  x"f6",  x"f0",  x"c3",  x"27",  x"f0", -- 1010
         x"c3",  x"7a",  x"f0",  x"c3",  x"99",  x"f0",  x"c5",  x"cd", -- 1018
         x"7a",  x"f0",  x"cd",  x"63",  x"f0",  x"18",  x"07",  x"c5", -- 1020
         x"cd",  x"7a",  x"f0",  x"cd",  x"77",  x"f0",  x"cd",  x"99", -- 1028
         x"f0",  x"c1",  x"c9",  x"f5",  x"db",  x"88",  x"cb",  x"d7", -- 1030
         x"d3",  x"88",  x"f1",  x"cd",  x"77",  x"f0",  x"f5",  x"db", -- 1038
         x"88",  x"cb",  x"97",  x"d3",  x"88",  x"f1",  x"c9",  x"f3", -- 1040
         x"e5",  x"e1",  x"e1",  x"23",  x"e5",  x"2b",  x"3b",  x"3b", -- 1048
         x"fb",  x"f5",  x"d5",  x"5e",  x"16",  x"00",  x"2a",  x"b0", -- 1050
         x"b7",  x"19",  x"19",  x"5e",  x"23",  x"56",  x"eb",  x"d1", -- 1058
         x"f1",  x"e3",  x"c9",  x"a7",  x"e5",  x"d5",  x"c5",  x"e5", -- 1060
         x"21",  x"bb",  x"f0",  x"e3",  x"e5",  x"f5",  x"d5",  x"38", -- 1068
         x"e3",  x"3a",  x"80",  x"b7",  x"5f",  x"18",  x"dd",  x"37", -- 1070
         x"18",  x"ea",  x"c1",  x"fd",  x"e5",  x"fd",  x"21",  x"00", -- 1078
         x"00",  x"fd",  x"39",  x"f3",  x"dd",  x"77",  x"0b",  x"db", -- 1080
         x"88",  x"cb",  x"d7",  x"cb",  x"ef",  x"d3",  x"88",  x"ed", -- 1088
         x"7b",  x"ae",  x"b7",  x"fb",  x"dd",  x"7e",  x"0b",  x"c5", -- 1090
         x"c9",  x"c1",  x"dd",  x"77",  x"0b",  x"db",  x"88",  x"cb", -- 1098
         x"97",  x"cb",  x"af",  x"f3",  x"d3",  x"88",  x"fd",  x"f9", -- 10A0
         x"fb",  x"dd",  x"7e",  x"0b",  x"fd",  x"e1",  x"c5",  x"c9", -- 10A8
         x"e3",  x"5e",  x"23",  x"56",  x"23",  x"eb",  x"19",  x"eb", -- 10B0
         x"e3",  x"d5",  x"c9",  x"c1",  x"d1",  x"e1",  x"c9",  x"31", -- 10B8
         x"c4",  x"01",  x"af",  x"47",  x"4f",  x"02",  x"0d",  x"20", -- 10C0
         x"fc",  x"10",  x"fa",  x"0e",  x"80",  x"ed",  x"79",  x"10", -- 10C8
         x"fc",  x"cd",  x"d0",  x"f3",  x"af",  x"32",  x"9b",  x"b7", -- 10D0
         x"cd",  x"bb",  x"f6",  x"3c",  x"fe",  x"0a",  x"38",  x"f5", -- 10D8
         x"cd",  x"8c",  x"f9",  x"3e",  x"0c",  x"cd",  x"29",  x"e3", -- 10E0
         x"cd",  x"6e",  x"f9",  x"cd",  x"61",  x"fb",  x"cd",  x"d9", -- 10E8
         x"c6",  x"cd",  x"6d",  x"fb",  x"18",  x"06",  x"31",  x"c4", -- 10F0
         x"01",  x"cd",  x"d0",  x"f3",  x"3a",  x"00",  x"a8",  x"3d", -- 10F8
         x"20",  x"0c",  x"cd",  x"61",  x"fb",  x"cd",  x"d5",  x"c2", -- 1100
         x"cd",  x"c3",  x"c6",  x"cd",  x"6d",  x"fb",  x"01",  x"80", -- 1108
         x"08",  x"ed",  x"78",  x"3d",  x"20",  x"1c",  x"3e",  x"43", -- 1110
         x"ed",  x"79",  x"32",  x"08",  x"b8",  x"dd",  x"7e",  x"04", -- 1118
         x"e6",  x"fc",  x"dd",  x"77",  x"04",  x"d3",  x"86",  x"c3", -- 1120
         x"00",  x"40",  x"7f",  x"7f",  x"4d",  x"45",  x"4e",  x"55", -- 1128
         x"01",  x"e1",  x"cd",  x"ee",  x"f1",  x"0c",  x"0a",  x"2a", -- 1130
         x"20",  x"4b",  x"43",  x"2d",  x"43",  x"41",  x"4f",  x"53", -- 1138
         x"20",  x"34",  x"2e",  x"32",  x"20",  x"2a",  x"00",  x"21", -- 1140
         x"00",  x"c0",  x"4d",  x"45",  x"cd",  x"6b",  x"f3",  x"cd", -- 1148
         x"ee",  x"f1",  x"02",  x"25",  x"00",  x"cd",  x"de",  x"e3", -- 1150
         x"38",  x"29",  x"dd",  x"7e",  x"09",  x"ed",  x"b1",  x"e2", -- 1158
         x"83",  x"f1",  x"ed",  x"a1",  x"20",  x"f7",  x"7e",  x"fe", -- 1160
         x"02",  x"38",  x"e1",  x"fe",  x"30",  x"38",  x"e0",  x"fe", -- 1168
         x"60",  x"30",  x"dc",  x"cd",  x"1d",  x"f2",  x"23",  x"0b", -- 1170
         x"18",  x"ec",  x"e1",  x"cd",  x"61",  x"f3",  x"cd",  x"ee", -- 1178
         x"f1",  x"25",  x"00",  x"cd",  x"34",  x"f3",  x"13",  x"1a", -- 1180
         x"fe",  x"20",  x"28",  x"f2",  x"a7",  x"28",  x"ef",  x"cd", -- 1188
         x"a9",  x"f1",  x"30",  x"e7",  x"e5",  x"cd",  x"c7",  x"f3", -- 1190
         x"38",  x"e0",  x"21",  x"7e",  x"f1",  x"e3",  x"7e",  x"23", -- 1198
         x"e5",  x"a7",  x"cd",  x"eb",  x"f4",  x"c0",  x"c3",  x"3e", -- 11A0
         x"f0",  x"21",  x"00",  x"c0",  x"45",  x"4d",  x"dd",  x"7e", -- 11A8
         x"09",  x"ed",  x"b1",  x"37",  x"3f",  x"e0",  x"ed",  x"a1", -- 11B0
         x"20",  x"f7",  x"f5",  x"d5",  x"1a",  x"13",  x"fe",  x"21", -- 11B8
         x"38",  x"08",  x"ed",  x"a1",  x"28",  x"f6",  x"d1",  x"f1", -- 11C0
         x"18",  x"e7",  x"7e",  x"fe",  x"02",  x"38",  x"07",  x"fe", -- 11C8
         x"20",  x"38",  x"f3",  x"23",  x"18",  x"f4",  x"f1",  x"f1", -- 11D0
         x"37",  x"c9",  x"3d",  x"c8",  x"f5",  x"f1",  x"18",  x"fa", -- 11D8
         x"47",  x"af",  x"cd",  x"da",  x"f1",  x"10",  x"fb",  x"c9", -- 11E0
         x"dd",  x"7e",  x"02",  x"cd",  x"76",  x"f3",  x"e3",  x"7e", -- 11E8
         x"23",  x"a7",  x"ca",  x"61",  x"f0",  x"cd",  x"1d",  x"f2", -- 11F0
         x"18",  x"f5",  x"cd",  x"0a",  x"f2",  x"21",  x"a0",  x"fb", -- 11F8
         x"e5",  x"2a",  x"b9",  x"b7",  x"e3",  x"22",  x"b9",  x"b7", -- 1200
         x"e1",  x"c9",  x"21",  x"a4",  x"fb",  x"e5",  x"2a",  x"bb", -- 1208
         x"b7",  x"e3",  x"22",  x"bb",  x"b7",  x"e1",  x"c9",  x"e5", -- 1210
         x"2a",  x"bb",  x"b7",  x"18",  x"04",  x"e5",  x"2a",  x"b9", -- 1218
         x"b7",  x"d5",  x"c5",  x"5e",  x"16",  x"00",  x"2a",  x"b0", -- 1220
         x"b7",  x"f5",  x"19",  x"19",  x"f1",  x"5e",  x"23",  x"56", -- 1228
         x"eb",  x"cd",  x"99",  x"e1",  x"c1",  x"d1",  x"e1",  x"c9", -- 1230
         x"e5",  x"d5",  x"c5",  x"dd",  x"cb",  x"08",  x"76",  x"20", -- 1238
         x"76",  x"ed",  x"5b",  x"a0",  x"b7",  x"cd",  x"6a",  x"e0", -- 1240
         x"af",  x"be",  x"28",  x"13",  x"5f",  x"cd",  x"4a",  x"f7", -- 1248
         x"1c",  x"06",  x"0f",  x"cd",  x"d5",  x"e3",  x"38",  x"1b", -- 1250
         x"0b",  x"78",  x"b1",  x"20",  x"f6",  x"18",  x"ee",  x"cd", -- 1258
         x"40",  x"e0",  x"cb",  x"cd",  x"cb",  x"d5",  x"7e",  x"47", -- 1260
         x"ee",  x"7f",  x"77",  x"cd",  x"d5",  x"e3",  x"30",  x"fb", -- 1268
         x"70",  x"18",  x"05",  x"cb",  x"43",  x"c4",  x"4a",  x"f7", -- 1270
         x"57",  x"dd",  x"cb",  x"08",  x"6e",  x"01",  x"07",  x"03", -- 1278
         x"c4",  x"05",  x"e3",  x"7a",  x"21",  x"a2",  x"b7",  x"cb", -- 1280
         x"66",  x"28",  x"0d",  x"ed",  x"5b",  x"a0",  x"b7",  x"cd", -- 1288
         x"63",  x"e1",  x"ed",  x"53",  x"a0",  x"b7",  x"18",  x"a9", -- 1290
         x"fe",  x"1b",  x"20",  x"04",  x"cb",  x"e6",  x"18",  x"a1", -- 1298
         x"fe",  x"f1",  x"38",  x"90",  x"dd",  x"cb",  x"08",  x"f6", -- 12A0
         x"e6",  x"0f",  x"47",  x"21",  x"00",  x"b9",  x"7e",  x"a7", -- 12A8
         x"23",  x"20",  x"fb",  x"10",  x"f9",  x"18",  x"08",  x"cd", -- 12B0
         x"de",  x"e3",  x"38",  x"1b",  x"2a",  x"d1",  x"b7",  x"7e", -- 12B8
         x"fe",  x"1b",  x"20",  x"0c",  x"23",  x"22",  x"d1",  x"b7", -- 12C0
         x"21",  x"a2",  x"b7",  x"cb",  x"e6",  x"c3",  x"3b",  x"f2", -- 12C8
         x"23",  x"22",  x"d1",  x"b7",  x"a7",  x"20",  x"07",  x"dd", -- 12D0
         x"cb",  x"08",  x"b6",  x"c3",  x"41",  x"f2",  x"21",  x"a2", -- 12D8
         x"b7",  x"cb",  x"66",  x"ca",  x"34",  x"f2",  x"ed",  x"5b", -- 12E0
         x"a0",  x"b7",  x"cd",  x"63",  x"e1",  x"ed",  x"53",  x"a0", -- 12E8
         x"b7",  x"c3",  x"3b",  x"f2",  x"22",  x"e3",  x"00",  x"00", -- 12F0
         x"00",  x"28",  x"20",  x"00",  x"00",  x"00",  x"39",  x"60", -- 12F8
         x"e2",  x"00",  x"ee",  x"00",  x"fe",  x"00",  x"ee",  x"00", -- 1300
         x"fe",  x"c4",  x"01",  x"a8",  x"fb",  x"c8",  x"fc",  x"d3", -- 1308
         x"88",  x"c3",  x"12",  x"f0",  x"a0",  x"fb",  x"a4",  x"fb", -- 1310
         x"c3",  x"53",  x"f3",  x"c3",  x"53",  x"f3",  x"c3",  x"53", -- 1318
         x"f3",  x"c3",  x"53",  x"f3",  x"82",  x"dc",  x"00",  x"b2", -- 1320
         x"db",  x"ed",  x"0b",  x"05",  x"00",  x"01",  x"a8",  x"08", -- 1328
         x"09",  x"a8",  x"09",  x"06",  x"cd",  x"17",  x"f2",  x"cd", -- 1330
         x"1d",  x"f2",  x"fe",  x"0d",  x"20",  x"f6",  x"cd",  x"6b", -- 1338
         x"f3",  x"ed",  x"5b",  x"a0",  x"b7",  x"ba",  x"20",  x"04", -- 1340
         x"3a",  x"9f",  x"b7",  x"57",  x"15",  x"e5",  x"cd",  x"6a", -- 1348
         x"e0",  x"eb",  x"e1",  x"c9",  x"7c",  x"cd",  x"76",  x"f3", -- 1350
         x"7d",  x"cd",  x"76",  x"f3",  x"3e",  x"20",  x"c3",  x"1d", -- 1358
         x"f2",  x"cd",  x"ee",  x"f1",  x"45",  x"52",  x"52",  x"4f", -- 1360
         x"52",  x"07",  x"00",  x"cd",  x"ee",  x"f1",  x"0d",  x"0a", -- 1368
         x"00",  x"c9",  x"3e",  x"10",  x"18",  x"e8",  x"f5",  x"1f", -- 1370
         x"1f",  x"1f",  x"1f",  x"cd",  x"7f",  x"f3",  x"f1",  x"e6", -- 1378
         x"0f",  x"c6",  x"90",  x"27",  x"ce",  x"40",  x"27",  x"18", -- 1380
         x"d5",  x"cd",  x"8c",  x"f3",  x"cd",  x"54",  x"f3",  x"eb", -- 1388
         x"c9",  x"13",  x"1a",  x"fe",  x"20",  x"28",  x"fa",  x"af", -- 1390
         x"21",  x"98",  x"b7",  x"77",  x"2b",  x"77",  x"2b",  x"77", -- 1398
         x"1a",  x"b7",  x"c8",  x"fe",  x"20",  x"c8",  x"d6",  x"30", -- 13A0
         x"d8",  x"fe",  x"0a",  x"38",  x"0b",  x"d6",  x"07",  x"e6", -- 13A8
         x"df",  x"fe",  x"0a",  x"d8",  x"fe",  x"10",  x"3f",  x"d8", -- 13B0
         x"13",  x"34",  x"23",  x"ed",  x"6f",  x"23",  x"ed",  x"6f", -- 13B8
         x"2b",  x"2b",  x"28",  x"dc",  x"1b",  x"37",  x"c9",  x"cd", -- 13C0
         x"61",  x"fb",  x"cd",  x"0e",  x"c7",  x"c3",  x"6d",  x"fb", -- 13C8
         x"11",  x"99",  x"b7",  x"21",  x"f4",  x"f2",  x"01",  x"34", -- 13D0
         x"00",  x"ed",  x"b0",  x"0e",  x"0c",  x"1e",  x"dd",  x"ed", -- 13D8
         x"b0",  x"21",  x"03",  x"01",  x"22",  x"00",  x"b8",  x"21", -- 13E0
         x"00",  x"03",  x"22",  x"02",  x"b8",  x"3e",  x"03",  x"32", -- 13E8
         x"04",  x"b8",  x"f3",  x"ed",  x"5e",  x"16",  x"07",  x"21", -- 13F0
         x"63",  x"f4",  x"cd",  x"5a",  x"f4",  x"dd",  x"21",  x"f0", -- 13F8
         x"01",  x"dd",  x"36",  x"01",  x"28",  x"dd",  x"36",  x"04", -- 1400
         x"63",  x"3e",  x"01",  x"21",  x"ba",  x"fc",  x"32",  x"d7", -- 1408
         x"b7",  x"1e",  x"e2",  x"57",  x"01",  x"0e",  x"00",  x"ed", -- 1410
         x"b0",  x"dd",  x"66",  x"01",  x"dd",  x"6e",  x"04",  x"d5", -- 1418
         x"dd",  x"e1",  x"dd",  x"36",  x"08",  x"88",  x"dd",  x"74", -- 1420
         x"01",  x"dd",  x"75",  x"04",  x"dd",  x"36",  x"0e",  x"3a", -- 1428
         x"dd",  x"36",  x"0f",  x"fc",  x"dd",  x"36",  x"09",  x"7f", -- 1430
         x"f3",  x"ed",  x"5e",  x"3a",  x"d7",  x"b7",  x"ed",  x"47", -- 1438
         x"16",  x"04",  x"21",  x"7b",  x"f4",  x"cd",  x"5a",  x"f4", -- 1440
         x"dd",  x"36",  x"05",  x"00",  x"dd",  x"36",  x"06",  x"b7", -- 1448
         x"c9",  x"c5",  x"4e",  x"23",  x"46",  x"23",  x"ed",  x"b3", -- 1450
         x"c1",  x"c9",  x"f3",  x"cd",  x"51",  x"f4",  x"15",  x"20", -- 1458
         x"fa",  x"fb",  x"c9",  x"8a",  x"01",  x"e4",  x"88",  x"01", -- 1460
         x"0f",  x"8a",  x"02",  x"0f",  x"03",  x"8b",  x"03",  x"e6", -- 1468
         x"0f",  x"83",  x"89",  x"01",  x"ff",  x"84",  x"01",  x"28", -- 1470
         x"86",  x"01",  x"63",  x"8a",  x"01",  x"e4",  x"8b",  x"01", -- 1478
         x"e6",  x"8c",  x"01",  x"e8",  x"8e",  x"02",  x"47",  x"0c", -- 1480
         x"7f",  x"7f",  x"53",  x"41",  x"56",  x"45",  x"01",  x"fe", -- 1488
         x"02",  x"da",  x"61",  x"f3",  x"cd",  x"ee",  x"f1",  x"4e", -- 1490
         x"41",  x"4d",  x"45",  x"20",  x"3a",  x"00",  x"cd",  x"34", -- 1498
         x"f3",  x"21",  x"06",  x"00",  x"19",  x"11",  x"00",  x"b7", -- 14A0
         x"01",  x"0b",  x"00",  x"ed",  x"b0",  x"af",  x"12",  x"21", -- 14A8
         x"81",  x"b7",  x"1e",  x"10",  x"0e",  x"15",  x"ed",  x"b0", -- 14B0
         x"cd",  x"48",  x"f4",  x"cd",  x"1c",  x"e5",  x"2a",  x"82", -- 14B8
         x"b7",  x"dd",  x"75",  x"05",  x"dd",  x"74",  x"06",  x"cd", -- 14C0
         x"ee",  x"f1",  x"02",  x"00",  x"cd",  x"e8",  x"f1",  x"00", -- 14C8
         x"01",  x"a0",  x"00",  x"cd",  x"de",  x"e3",  x"da",  x"e0", -- 14D0
         x"e4",  x"11",  x"80",  x"00",  x"19",  x"ed",  x"5b",  x"84", -- 14D8
         x"b7",  x"ed",  x"52",  x"d2",  x"d9",  x"e4",  x"cd",  x"2b", -- 14E0
         x"e5",  x"18",  x"d6",  x"ed",  x"4b",  x"86",  x"b7",  x"ed", -- 14E8
         x"5b",  x"84",  x"b7",  x"2a",  x"82",  x"b7",  x"3a",  x"81", -- 14F0
         x"b7",  x"c9",  x"dd",  x"34",  x"03",  x"cd",  x"91",  x"e5", -- 14F8
         x"30",  x"20",  x"cd",  x"ee",  x"f1",  x"09",  x"09",  x"09", -- 1500
         x"20",  x"00",  x"cd",  x"e8",  x"f1",  x"20",  x"3f",  x"1e", -- 1508
         x"00",  x"dd",  x"7e",  x"03",  x"3d",  x"28",  x"e6",  x"cd", -- 1510
         x"38",  x"f2",  x"fe",  x"03",  x"37",  x"c8",  x"fe",  x"0a", -- 1518
         x"20",  x"db",  x"dd",  x"7e",  x"02",  x"dd",  x"46",  x"03", -- 1520
         x"05",  x"28",  x"17",  x"04",  x"b8",  x"28",  x"0b",  x"3c", -- 1528
         x"28",  x"08",  x"cd",  x"e8",  x"f1",  x"2a",  x"19",  x"00", -- 1530
         x"18",  x"c3",  x"cd",  x"e8",  x"f1",  x"3e",  x"20",  x"19", -- 1538
         x"00",  x"c9",  x"3d",  x"20",  x"ed",  x"cd",  x"6b",  x"f3", -- 1540
         x"21",  x"00",  x"b7",  x"06",  x"0b",  x"7e",  x"23",  x"cd", -- 1548
         x"29",  x"e3",  x"10",  x"f9",  x"c3",  x"5c",  x"f3",  x"cd", -- 1550
         x"ee",  x"f1",  x"3f",  x"3f",  x"3f",  x"00",  x"c3",  x"e0", -- 1558
         x"e4",  x"7f",  x"7f",  x"56",  x"45",  x"52",  x"49",  x"46", -- 1560
         x"59",  x"01",  x"dd",  x"cb",  x"07",  x"86",  x"18",  x"0b", -- 1568
         x"7f",  x"7f",  x"4c",  x"4f",  x"41",  x"44",  x"01",  x"dd", -- 1570
         x"cb",  x"07",  x"c6",  x"cd",  x"b4",  x"e4",  x"cd",  x"48", -- 1578
         x"f4",  x"dd",  x"36",  x"03",  x"00",  x"cd",  x"fa",  x"f4", -- 1580
         x"38",  x"d4",  x"dd",  x"cb",  x"07",  x"46",  x"28",  x"49", -- 1588
         x"2e",  x"10",  x"dd",  x"7e",  x"07",  x"e6",  x"e3",  x"dd", -- 1590
         x"77",  x"07",  x"7e",  x"cb",  x"27",  x"cb",  x"27",  x"e6", -- 1598
         x"1c",  x"dd",  x"b6",  x"07",  x"dd",  x"77",  x"07",  x"7e", -- 15A0
         x"d6",  x"02",  x"fe",  x"09",  x"30",  x"a9",  x"ed",  x"4b", -- 15A8
         x"15",  x"b7",  x"ed",  x"5b",  x"13",  x"b7",  x"2a",  x"11", -- 15B0
         x"b7",  x"3a",  x"81",  x"b7",  x"a7",  x"28",  x"13",  x"c5", -- 15B8
         x"ed",  x"4b",  x"82",  x"b7",  x"09",  x"eb",  x"09",  x"eb", -- 15C0
         x"dd",  x"cb",  x"07",  x"66",  x"20",  x"03",  x"e3",  x"09", -- 15C8
         x"e3",  x"c1",  x"ed",  x"43",  x"84",  x"b7",  x"cd",  x"89", -- 15D0
         x"f3",  x"cd",  x"6b",  x"f3",  x"eb",  x"cd",  x"fa",  x"f4", -- 15D8
         x"38",  x"a6",  x"dd",  x"cb",  x"07",  x"46",  x"28",  x"12", -- 15E0
         x"e5",  x"ed",  x"52",  x"01",  x"80",  x"00",  x"ed",  x"42", -- 15E8
         x"09",  x"30",  x"01",  x"4d",  x"21",  x"00",  x"b7",  x"ed", -- 15F0
         x"b0",  x"e1",  x"dd",  x"34",  x"02",  x"20",  x"de",  x"cd", -- 15F8
         x"e0",  x"e4",  x"dd",  x"7e",  x"07",  x"e6",  x"03",  x"3d", -- 1600
         x"c0",  x"dd",  x"7e",  x"07",  x"e6",  x"1c",  x"fe",  x"0c", -- 1608
         x"dd",  x"36",  x"07",  x"00",  x"d8",  x"2a",  x"84",  x"b7", -- 1610
         x"e9",  x"7f",  x"7f",  x"43",  x"4f",  x"4c",  x"4f",  x"52", -- 1618
         x"01",  x"cd",  x"61",  x"fb",  x"cd",  x"63",  x"c1",  x"c3", -- 1620
         x"6d",  x"fb",  x"e5",  x"21",  x"a2",  x"b7",  x"cb",  x"de", -- 1628
         x"cd",  x"1d",  x"f2",  x"cb",  x"9e",  x"e1",  x"c9",  x"7f", -- 1630
         x"7f",  x"44",  x"49",  x"53",  x"50",  x"4c",  x"41",  x"59", -- 1638
         x"01",  x"cd",  x"61",  x"fb",  x"cd",  x"42",  x"c2",  x"c3", -- 1640
         x"6d",  x"fb",  x"cd",  x"6d",  x"fb",  x"7e",  x"c3",  x"61", -- 1648
         x"fb",  x"7f",  x"7f",  x"4d",  x"4f",  x"44",  x"49",  x"46", -- 1650
         x"59",  x"01",  x"cd",  x"61",  x"fb",  x"cd",  x"6a",  x"c2", -- 1658
         x"18",  x"e5",  x"cd",  x"6d",  x"fb",  x"77",  x"18",  x"e6", -- 1660
         x"7f",  x"7f",  x"57",  x"49",  x"4e",  x"44",  x"4f",  x"57", -- 1668
         x"01",  x"a7",  x"28",  x"2a",  x"3d",  x"28",  x"26",  x"65", -- 1670
         x"69",  x"53",  x"3a",  x"88",  x"b7",  x"5f",  x"3a",  x"81", -- 1678
         x"b7",  x"fe",  x"04",  x"20",  x"05",  x"38",  x"09",  x"af", -- 1680
         x"18",  x"03",  x"3a",  x"8a",  x"b7",  x"cd",  x"94",  x"f6", -- 1688
         x"da",  x"61",  x"f3",  x"c9",  x"cd",  x"61",  x"fb",  x"cd", -- 1690
         x"2d",  x"c1",  x"c3",  x"6d",  x"fb",  x"7d",  x"cd",  x"bb", -- 1698
         x"f6",  x"32",  x"9b",  x"b7",  x"cd",  x"ae",  x"f6",  x"d8", -- 16A0
         x"eb",  x"11",  x"9c",  x"b7",  x"18",  x"1b",  x"c6",  x"f6", -- 16A8
         x"d8",  x"87",  x"5f",  x"87",  x"87",  x"83",  x"5f",  x"16", -- 16B0
         x"b9",  x"a7",  x"c9",  x"f5",  x"3a",  x"9b",  x"b7",  x"cd", -- 16B8
         x"ae",  x"f6",  x"da",  x"5b",  x"e0",  x"f1",  x"21",  x"9c", -- 16C0
         x"b7",  x"01",  x"0a",  x"00",  x"ed",  x"b0",  x"c9",  x"23", -- 16C8
         x"7e",  x"a7",  x"c8",  x"cd",  x"2a",  x"f6",  x"18",  x"f7", -- 16D0
         x"7f",  x"7f",  x"4b",  x"45",  x"59",  x"01",  x"fe",  x"01", -- 16D8
         x"c0",  x"7d",  x"a7",  x"c8",  x"fe",  x"0d",  x"d0",  x"47", -- 16E0
         x"21",  x"00",  x"b9",  x"7e",  x"23",  x"a7",  x"20",  x"fb", -- 16E8
         x"10",  x"f9",  x"cd",  x"d0",  x"f6",  x"f5",  x"2b",  x"f1", -- 16F0
         x"cd",  x"17",  x"f2",  x"fe",  x"13",  x"ca",  x"6b",  x"f3", -- 16F8
         x"f5",  x"06",  x"00",  x"3d",  x"20",  x"15",  x"7e",  x"a7", -- 1700
         x"28",  x"ed",  x"54",  x"5d",  x"e5",  x"23",  x"3e",  x"9c", -- 1708
         x"95",  x"4f",  x"ed",  x"b0",  x"e1",  x"f1",  x"cd",  x"1d", -- 1710
         x"f2",  x"18",  x"da",  x"3a",  x"9a",  x"b9",  x"a7",  x"20", -- 1718
         x"d6",  x"e5",  x"3e",  x"9b",  x"95",  x"4f",  x"21",  x"9a", -- 1720
         x"b9",  x"11",  x"9b",  x"b9",  x"ed",  x"b8",  x"e1",  x"f1", -- 1728
         x"23",  x"77",  x"cd",  x"2a",  x"f6",  x"18",  x"c1",  x"7f", -- 1730
         x"7f",  x"4b",  x"45",  x"59",  x"4c",  x"49",  x"53",  x"54", -- 1738
         x"01",  x"cd",  x"61",  x"fb",  x"cd",  x"f7",  x"c0",  x"c3", -- 1740
         x"6d",  x"fb",  x"d5",  x"f5",  x"e5",  x"cd",  x"40",  x"e0", -- 1748
         x"38",  x"0a",  x"c5",  x"06",  x"08",  x"7e",  x"2f",  x"77", -- 1750
         x"2c",  x"10",  x"fa",  x"c1",  x"e1",  x"f1",  x"d1",  x"c9", -- 1758
         x"e5",  x"d5",  x"c5",  x"a7",  x"f5",  x"2a",  x"d3",  x"b7", -- 1760
         x"ed",  x"5b",  x"d5",  x"b7",  x"16",  x"00",  x"c3",  x"ec", -- 1768
         x"f7",  x"cd",  x"61",  x"fb",  x"cd",  x"e4",  x"c1",  x"c3", -- 1770
         x"6d",  x"fb",  x"3a",  x"86",  x"b7",  x"4f",  x"69",  x"af", -- 1778
         x"06",  x"08",  x"cb",  x"1d",  x"30",  x"01",  x"81",  x"1f", -- 1780
         x"cb",  x"1d",  x"10",  x"f8",  x"67",  x"54",  x"5d",  x"79", -- 1788
         x"cb",  x"21",  x"cb",  x"10",  x"0b",  x"c5",  x"01",  x"01", -- 1790
         x"00",  x"d9",  x"4f",  x"06",  x"00",  x"cd",  x"c2",  x"f7", -- 1798
         x"cd",  x"c2",  x"f7",  x"d9",  x"a7",  x"ed",  x"42",  x"03", -- 17A0
         x"03",  x"ed",  x"52",  x"19",  x"d9",  x"30",  x"0c",  x"d9", -- 17A8
         x"e3",  x"eb",  x"a7",  x"ed",  x"52",  x"1b",  x"1b",  x"eb", -- 17B0
         x"e3",  x"d9",  x"0d",  x"04",  x"79",  x"b8",  x"30",  x"dd", -- 17B8
         x"f1",  x"c9",  x"78",  x"41",  x"4f",  x"af",  x"57",  x"2a", -- 17C0
         x"84",  x"b7",  x"e5",  x"59",  x"19",  x"cd",  x"d6",  x"f7", -- 17C8
         x"af",  x"57",  x"e1",  x"59",  x"ed",  x"52",  x"e5",  x"2a", -- 17D0
         x"82",  x"b7",  x"58",  x"a7",  x"ed",  x"52",  x"d1",  x"cd", -- 17D8
         x"e8",  x"f7",  x"d5",  x"57",  x"58",  x"19",  x"19",  x"d1", -- 17E0
         x"e5",  x"d5",  x"c5",  x"f5",  x"7d",  x"e6",  x"07",  x"c6", -- 17E8
         x"f8",  x"4f",  x"06",  x"fd",  x"7d",  x"cb",  x"3c",  x"1f", -- 17F0
         x"cb",  x"3c",  x"1f",  x"cb",  x"3c",  x"1f",  x"fe",  x"28", -- 17F8
         x"30",  x"31",  x"f6",  x"80",  x"67",  x"3e",  x"ff",  x"82", -- 1800
         x"38",  x"29",  x"ab",  x"6f",  x"3a",  x"d6",  x"b7",  x"57", -- 1808
         x"0a",  x"dd",  x"cb",  x"01",  x"5e",  x"28",  x"2d",  x"cb", -- 1810
         x"4a",  x"20",  x"23",  x"cb",  x"42",  x"20",  x"19",  x"b6", -- 1818
         x"77",  x"dd",  x"7e",  x"01",  x"5f",  x"ee",  x"02",  x"f3", -- 1820
         x"d3",  x"84",  x"7e",  x"e6",  x"07",  x"b2",  x"77",  x"7b", -- 1828
         x"d3",  x"84",  x"fb",  x"f1",  x"c1",  x"d1",  x"e1",  x"c9", -- 1830
         x"ae",  x"cb",  x"82",  x"c3",  x"20",  x"f8",  x"2f",  x"a6", -- 1838
         x"77",  x"c3",  x"33",  x"f8",  x"47",  x"b6",  x"cb",  x"5a", -- 1840
         x"20",  x"01",  x"a8",  x"77",  x"dd",  x"7e",  x"01",  x"4f", -- 1848
         x"ee",  x"02",  x"f3",  x"d3",  x"84",  x"78",  x"b6",  x"cb", -- 1850
         x"62",  x"20",  x"01",  x"a8",  x"77",  x"79",  x"d3",  x"84", -- 1858
         x"fb",  x"18",  x"d0",  x"cd",  x"61",  x"fb",  x"cd",  x"7c", -- 1860
         x"c1",  x"18",  x"28",  x"cd",  x"61",  x"fb",  x"cd",  x"2b", -- 1868
         x"c7",  x"18",  x"20",  x"cd",  x"61",  x"fb",  x"cd",  x"a7", -- 1870
         x"c7",  x"18",  x"18",  x"cd",  x"6d",  x"fb",  x"2a",  x"c9", -- 1878
         x"b7",  x"cd",  x"99",  x"f0",  x"e9",  x"7f",  x"7f",  x"4d", -- 1880
         x"4f",  x"44",  x"55",  x"4c",  x"01",  x"cd",  x"61",  x"fb", -- 1888
         x"cd",  x"00",  x"c0",  x"c3",  x"6d",  x"fb",  x"7f",  x"7f", -- 1890
         x"53",  x"59",  x"53",  x"54",  x"45",  x"4d",  x"01",  x"cd", -- 1898
         x"61",  x"fb",  x"cd",  x"28",  x"c0",  x"18",  x"ec",  x"e5", -- 18A0
         x"c5",  x"cd",  x"7a",  x"f0",  x"cb",  x"6b",  x"d5",  x"20", -- 18A8
         x"53",  x"23",  x"23",  x"cb",  x"7b",  x"20",  x"42",  x"e5", -- 18B0
         x"7b",  x"e6",  x"07",  x"21",  x"f1",  x"f8",  x"85",  x"6f", -- 18B8
         x"7a",  x"53",  x"5e",  x"e1",  x"cd",  x"77",  x"f0",  x"d1", -- 18C0
         x"57",  x"7b",  x"e6",  x"4f",  x"ee",  x"43",  x"20",  x"18", -- 18C8
         x"cd",  x"ee",  x"f1",  x"56",  x"45",  x"52",  x"49",  x"46", -- 18D0
         x"59",  x"20",  x"3f",  x"28",  x"59",  x"29",  x"3a",  x"00", -- 18D8
         x"cd",  x"38",  x"f2",  x"fe",  x"59",  x"cc",  x"6a",  x"f5", -- 18E0
         x"7a",  x"cb",  x"9b",  x"cd",  x"99",  x"f0",  x"c1",  x"e1", -- 18E8
         x"c9",  x"16",  x"24",  x"37",  x"38",  x"06",  x"02",  x"07", -- 18F0
         x"03",  x"cd",  x"ca",  x"e3",  x"d1",  x"57",  x"30",  x"e8", -- 18F8
         x"cb",  x"bb",  x"18",  x"e4",  x"3a",  x"5e",  x"03",  x"a7", -- 1900
         x"28",  x"09",  x"cd",  x"99",  x"f0",  x"cd",  x"41",  x"c6", -- 1908
         x"cd",  x"7a",  x"f0",  x"db",  x"88",  x"e6",  x"5f",  x"d3", -- 1910
         x"88",  x"c3",  x"7e",  x"f1",  x"7e",  x"23",  x"a7",  x"c8", -- 1918
         x"cd",  x"1d",  x"f2",  x"18",  x"f7",  x"cd",  x"eb",  x"f4", -- 1920
         x"dd",  x"cb",  x"08",  x"4e",  x"20",  x"fa",  x"c5",  x"0e", -- 1928
         x"8c",  x"cd",  x"5a",  x"f9",  x"0c",  x"eb",  x"cd",  x"5a", -- 1930
         x"f9",  x"c1",  x"79",  x"ee",  x"1f",  x"f6",  x"81",  x"4f", -- 1938
         x"78",  x"a7",  x"28",  x"0d",  x"cb",  x"b9",  x"dd",  x"cb", -- 1940
         x"08",  x"ce",  x"3e",  x"c7",  x"d3",  x"8e",  x"78",  x"d3", -- 1948
         x"8e",  x"06",  x"60",  x"db",  x"89",  x"a0",  x"b1",  x"d3", -- 1950
         x"89",  x"c9",  x"7d",  x"a7",  x"2e",  x"03",  x"28",  x"0b", -- 1958
         x"6f",  x"3e",  x"07",  x"cb",  x"44",  x"28",  x"02",  x"f6", -- 1960
         x"20",  x"ed",  x"79",  x"ed",  x"69",  x"c9",  x"21",  x"00", -- 1968
         x"b2",  x"22",  x"cb",  x"b7",  x"dd",  x"7e",  x"01",  x"e6", -- 1970
         x"f8",  x"d3",  x"84",  x"dd",  x"77",  x"01",  x"c9",  x"21", -- 1978
         x"00",  x"ad",  x"22",  x"cb",  x"b7",  x"dd",  x"7e",  x"01", -- 1980
         x"f6",  x"05",  x"18",  x"ed",  x"21",  x"00",  x"ad",  x"22", -- 1988
         x"cb",  x"b7",  x"dd",  x"7e",  x"01",  x"e6",  x"fe",  x"f6", -- 1990
         x"04",  x"18",  x"de",  x"21",  x"00",  x"b2",  x"22",  x"cb", -- 1998
         x"b7",  x"dd",  x"7e",  x"01",  x"f6",  x"01",  x"e6",  x"f9", -- 19A0
         x"18",  x"cf",  x"21",  x"a2",  x"b7",  x"7e",  x"ee",  x"04", -- 19A8
         x"77",  x"c9",  x"dd",  x"7e",  x"01",  x"ee",  x"02",  x"18", -- 19B0
         x"c0",  x"db",  x"89",  x"ee",  x"80",  x"d3",  x"89",  x"dd", -- 19B8
         x"7e",  x"01",  x"ee",  x"08",  x"18",  x"b3",  x"7f",  x"7f", -- 19C0
         x"56",  x"32",  x"34",  x"4f",  x"55",  x"54",  x"01",  x"cd", -- 19C8
         x"61",  x"fb",  x"cd",  x"d5",  x"c2",  x"3e",  x"0d",  x"cd", -- 19D0
         x"06",  x"fa",  x"3e",  x"0a",  x"cd",  x"06",  x"fa",  x"c3", -- 19D8
         x"6d",  x"fb",  x"cd",  x"61",  x"fb",  x"cd",  x"cf",  x"c3", -- 19E0
         x"18",  x"f5",  x"7f",  x"7f",  x"56",  x"32",  x"34",  x"44", -- 19E8
         x"55",  x"50",  x"01",  x"cd",  x"61",  x"fb",  x"cd",  x"4f", -- 19F0
         x"c6",  x"18",  x"e4",  x"cd",  x"61",  x"fb",  x"cd",  x"c3", -- 19F8
         x"c6",  x"18",  x"dc",  x"cd",  x"29",  x"e3",  x"f5",  x"3a", -- 1A00
         x"e1",  x"b7",  x"cb",  x"7f",  x"28",  x"29",  x"e6",  x"f0", -- 1A08
         x"fe",  x"90",  x"28",  x"17",  x"fe",  x"a0",  x"20",  x"1f", -- 1A10
         x"f1",  x"e5",  x"c5",  x"21",  x"92",  x"fb",  x"01",  x"07", -- 1A18
         x"00",  x"ed",  x"b1",  x"20",  x"0f",  x"0e",  x"06",  x"09", -- 1A20
         x"7e",  x"18",  x"09",  x"f1",  x"fe",  x"7e",  x"20",  x"08", -- 1A28
         x"3e",  x"83",  x"18",  x"04",  x"c1",  x"e1",  x"f5",  x"f1", -- 1A30
         x"fe",  x"09",  x"28",  x"0d",  x"f5",  x"3a",  x"a2",  x"b7", -- 1A38
         x"cb",  x"5f",  x"28",  x"0e",  x"f1",  x"fe",  x"7f",  x"20", -- 1A40
         x"02",  x"3e",  x"20",  x"fe",  x"20",  x"30",  x"02",  x"3e", -- 1A48
         x"5f",  x"f5",  x"c5",  x"cd",  x"d4",  x"fa",  x"3e",  x"0a", -- 1A50
         x"81",  x"4f",  x"ed",  x"78",  x"cb",  x"57",  x"20",  x"08", -- 1A58
         x"3e",  x"01",  x"cd",  x"e0",  x"f1",  x"c1",  x"18",  x"ea", -- 1A60
         x"c1",  x"f1",  x"c5",  x"f5",  x"cd",  x"d4",  x"fa",  x"3e", -- 1A68
         x"08",  x"81",  x"4f",  x"f1",  x"ed",  x"79",  x"c1",  x"c9", -- 1A70
         x"f5",  x"c5",  x"cd",  x"e1",  x"fa",  x"3e",  x"0a",  x"81", -- 1A78
         x"4f",  x"ed",  x"78",  x"cb",  x"57",  x"20",  x"08",  x"3e", -- 1A80
         x"01",  x"cd",  x"e0",  x"f1",  x"c1",  x"18",  x"ea",  x"c1", -- 1A88
         x"f1",  x"c5",  x"f5",  x"cd",  x"e1",  x"fa",  x"18",  x"d7", -- 1A90
         x"c5",  x"e5",  x"d5",  x"cd",  x"e1",  x"fa",  x"c5",  x"3e", -- 1A98
         x"0a",  x"81",  x"4f",  x"ed",  x"78",  x"cb",  x"47",  x"20", -- 1AA0
         x"15",  x"3e",  x"05",  x"ed",  x"79",  x"3e",  x"ea",  x"ed", -- 1AA8
         x"79",  x"ed",  x"78",  x"cb",  x"47",  x"20",  x"07",  x"cd", -- 1AB0
         x"de",  x"e3",  x"38",  x"15",  x"18",  x"f3",  x"3e",  x"05", -- 1AB8
         x"ed",  x"79",  x"3e",  x"6a",  x"ed",  x"79",  x"c1",  x"3e", -- 1AC0
         x"08",  x"81",  x"4f",  x"ed",  x"78",  x"d1",  x"e1",  x"c1", -- 1AC8
         x"c9",  x"c1",  x"18",  x"f9",  x"f5",  x"3a",  x"e1",  x"b7", -- 1AD0
         x"cb",  x"57",  x"0e",  x"01",  x"20",  x"01",  x"0d",  x"f1", -- 1AD8
         x"c9",  x"f5",  x"3a",  x"e8",  x"b7",  x"18",  x"f1",  x"e5", -- 1AE0
         x"d5",  x"c5",  x"f5",  x"db",  x"09",  x"f5",  x"3e",  x"18", -- 1AE8
         x"d3",  x"0b",  x"3e",  x"05",  x"d3",  x"0b",  x"3e",  x"6a", -- 1AF0
         x"d3",  x"0b",  x"f1",  x"cd",  x"57",  x"fb",  x"fe",  x"0d", -- 1AF8
         x"28",  x"0a",  x"fe",  x"1b",  x"28",  x"13",  x"cd",  x"fb", -- 1B00
         x"f9",  x"c3",  x"24",  x"e1",  x"cd",  x"fb",  x"f9",  x"21", -- 1B08
         x"5a",  x"fb",  x"f3",  x"22",  x"e2",  x"01",  x"fb",  x"18", -- 1B10
         x"f0",  x"3e",  x"06",  x"32",  x"e8",  x"b7",  x"cd",  x"f3", -- 1B18
         x"f9",  x"cd",  x"98",  x"fa",  x"fe",  x"54",  x"28",  x"06", -- 1B20
         x"fe",  x"55",  x"28",  x"1e",  x"18",  x"d8",  x"cd",  x"98", -- 1B28
         x"fa",  x"6f",  x"cd",  x"98",  x"fa",  x"67",  x"cd",  x"98", -- 1B30
         x"fa",  x"4f",  x"cd",  x"98",  x"fa",  x"47",  x"cd",  x"98", -- 1B38
         x"fa",  x"77",  x"23",  x"0b",  x"79",  x"b0",  x"20",  x"f6", -- 1B40
         x"18",  x"bc",  x"cd",  x"98",  x"fa",  x"6f",  x"cd",  x"98", -- 1B48
         x"fa",  x"67",  x"cd",  x"99",  x"e1",  x"18",  x"af",  x"fb", -- 1B50
         x"ed",  x"4d",  x"fb",  x"f5",  x"db",  x"09",  x"c3",  x"b5", -- 1B58
         x"e3",  x"f5",  x"dd",  x"cb",  x"04",  x"fe",  x"dd",  x"7e", -- 1B60
         x"04",  x"d3",  x"86",  x"f1",  x"c9",  x"f5",  x"dd",  x"cb", -- 1B68
         x"04",  x"be",  x"dd",  x"7e",  x"04",  x"d3",  x"86",  x"f1", -- 1B70
         x"c9",  x"cd",  x"61",  x"fb",  x"cd",  x"1c",  x"c1",  x"18", -- 1B78
         x"ec",  x"cd",  x"61",  x"fb",  x"cd",  x"0e",  x"c1",  x"18", -- 1B80
         x"e4",  x"cd",  x"17",  x"e6",  x"f5",  x"cd",  x"cd",  x"e4", -- 1B88
         x"f1",  x"c9",  x"7b",  x"7c",  x"7d",  x"7e",  x"5b",  x"5c", -- 1B90
         x"5d",  x"84",  x"94",  x"81",  x"e1",  x"8e",  x"99",  x"9a", -- 1B98
         x"00",  x"38",  x"02",  x"03",  x"04",  x"37",  x"06",  x"07", -- 1BA0
         x"29",  x"e3",  x"2b",  x"e5",  x"bd",  x"b7",  x"c3",  x"b7", -- 1BA8
         x"38",  x"f2",  x"91",  x"e5",  x"c0",  x"b7",  x"c6",  x"b7", -- 1BB0
         x"1c",  x"e5",  x"d9",  x"e4",  x"8e",  x"e5",  x"ff",  x"f5", -- 1BB8
         x"ca",  x"e3",  x"f6",  x"f0",  x"d5",  x"e3",  x"21",  x"f6", -- 1BC0
         x"77",  x"f5",  x"6a",  x"f5",  x"7e",  x"f1",  x"fa",  x"f1", -- 1BC8
         x"e0",  x"f1",  x"eb",  x"f4",  x"17",  x"f2",  x"34",  x"f3", -- 1BD0
         x"92",  x"f3",  x"61",  x"f3",  x"54",  x"f3",  x"89",  x"f3", -- 1BD8
         x"76",  x"f3",  x"b1",  x"f1",  x"00",  x"f2",  x"0d",  x"f2", -- 1BE0
         x"fd",  x"f1",  x"0a",  x"f2",  x"c7",  x"f3",  x"ee",  x"f1", -- 1BE8
         x"1d",  x"f2",  x"4a",  x"f7",  x"04",  x"e4",  x"9b",  x"e4", -- 1BF0
         x"16",  x"e3",  x"18",  x"e3",  x"de",  x"e3",  x"5c",  x"f3", -- 1BF8
         x"6b",  x"f3",  x"72",  x"f3",  x"5a",  x"f6",  x"71",  x"f7", -- 1C00
         x"60",  x"f7",  x"0b",  x"f4",  x"6a",  x"e0",  x"5e",  x"e0", -- 1C08
         x"4e",  x"e0",  x"25",  x"f9",  x"a5",  x"f4",  x"73",  x"f8", -- 1C10
         x"6b",  x"f8",  x"e2",  x"f6",  x"41",  x"f7",  x"41",  x"f6", -- 1C18
         x"94",  x"f6",  x"9e",  x"f6",  x"63",  x"f8",  x"7a",  x"f7", -- 1C20
         x"81",  x"fb",  x"79",  x"fb",  x"2a",  x"f6",  x"51",  x"f4", -- 1C28
         x"5a",  x"f4",  x"1c",  x"f9",  x"47",  x"f1",  x"cf",  x"f9", -- 1C30
         x"f3",  x"f9",  x"57",  x"77",  x"41",  x"61",  x"32",  x"22", -- 1C38
         x"08",  x"19",  x"10",  x"0c",  x"2d",  x"3d",  x"f2",  x"f8", -- 1C40
         x"59",  x"79",  x"45",  x"65",  x"53",  x"73",  x"33",  x"23", -- 1C48
         x"5e",  x"5d",  x"01",  x"0f",  x"3a",  x"2a",  x"f3",  x"f9", -- 1C50
         x"58",  x"78",  x"54",  x"74",  x"46",  x"66",  x"35",  x"25", -- 1C58
         x"50",  x"70",  x"1f",  x"02",  x"30",  x"40",  x"f5",  x"fb", -- 1C60
         x"56",  x"76",  x"55",  x"75",  x"48",  x"68",  x"37",  x"27", -- 1C68
         x"4f",  x"6f",  x"1a",  x"14",  x"39",  x"29",  x"03",  x"03", -- 1C70
         x"4e",  x"6e",  x"49",  x"69",  x"4a",  x"6a",  x"38",  x"28", -- 1C78
         x"20",  x"5b",  x"4b",  x"6b",  x"2c",  x"3c",  x"13",  x"1b", -- 1C80
         x"4d",  x"6d",  x"5a",  x"7a",  x"47",  x"67",  x"36",  x"26", -- 1C88
         x"00",  x"00",  x"4c",  x"6c",  x"2e",  x"3e",  x"f6",  x"fc", -- 1C90
         x"42",  x"62",  x"52",  x"72",  x"44",  x"64",  x"34",  x"24", -- 1C98
         x"5f",  x"5c",  x"2b",  x"3b",  x"2f",  x"3f",  x"f4",  x"fa", -- 1CA0
         x"43",  x"63",  x"51",  x"71",  x"16",  x"16",  x"31",  x"21", -- 1CA8
         x"0a",  x"12",  x"0b",  x"11",  x"09",  x"18",  x"f1",  x"f7", -- 1CB0
         x"0d",  x"0d",  x"e7",  x"fa",  x"08",  x"e6",  x"45",  x"e3", -- 1CB8
         x"17",  x"e6",  x"f8",  x"e5",  x"89",  x"fb",  x"39",  x"e3", -- 1CC0
         x"22",  x"e3",  x"e2",  x"e1",  x"aa",  x"e2",  x"22",  x"e3", -- 1CC8
         x"22",  x"e3",  x"22",  x"e3",  x"22",  x"e3",  x"eb",  x"e2", -- 1CD0
         x"c1",  x"e1",  x"aa",  x"e1",  x"b3",  x"e1",  x"d1",  x"e1", -- 1CD8
         x"37",  x"e2",  x"47",  x"e2",  x"22",  x"e3",  x"bd",  x"e1", -- 1CE0
         x"45",  x"e2",  x"d6",  x"e1",  x"dd",  x"e1",  x"22",  x"e3", -- 1CE8
         x"1a",  x"e3",  x"22",  x"e3",  x"22",  x"e3",  x"22",  x"e3", -- 1CF0
         x"cb",  x"e1",  x"47",  x"e2",  x"18",  x"e2",  x"23",  x"e3", -- 1CF8
         x"22",  x"e3",  x"22",  x"e3",  x"b1",  x"e1",  x"e5",  x"e1", -- 1D00
         x"c9",  x"4e",  x"4b",  x"45",  x"59",  x"24",  x"ca",  x"4f", -- 1D08
         x"59",  x"53",  x"54",  x"d3",  x"54",  x"52",  x"49",  x"4e", -- 1D10
         x"47",  x"24",  x"c9",  x"4e",  x"53",  x"54",  x"52",  x"d2", -- 1D18
         x"45",  x"4e",  x"55",  x"4d",  x"42",  x"45",  x"52",  x"c4", -- 1D20
         x"45",  x"4c",  x"45",  x"54",  x"45",  x"d0",  x"41",  x"55", -- 1D28
         x"53",  x"45",  x"c2",  x"45",  x"45",  x"50",  x"d7",  x"49", -- 1D30
         x"4e",  x"44",  x"4f",  x"57",  x"c2",  x"4f",  x"52",  x"44", -- 1D38
         x"45",  x"52",  x"c9",  x"4e",  x"4b",  x"d0",  x"41",  x"50", -- 1D40
         x"45",  x"52",  x"c1",  x"54",  x"c3",  x"4f",  x"4c",  x"4f", -- 1D48
         x"52",  x"d3",  x"4f",  x"55",  x"4e",  x"44",  x"d0",  x"53", -- 1D50
         x"45",  x"54",  x"d0",  x"52",  x"45",  x"53",  x"45",  x"54", -- 1D58
         x"c2",  x"4c",  x"4f",  x"41",  x"44",  x"d6",  x"50",  x"45", -- 1D60
         x"45",  x"4b",  x"d6",  x"50",  x"4f",  x"4b",  x"45",  x"cc", -- 1D68
         x"4f",  x"43",  x"41",  x"54",  x"45",  x"cb",  x"45",  x"59", -- 1D70
         x"4c",  x"49",  x"53",  x"54",  x"cb",  x"45",  x"59",  x"d3", -- 1D78
         x"57",  x"49",  x"54",  x"43",  x"48",  x"d0",  x"54",  x"45", -- 1D80
         x"53",  x"54",  x"c3",  x"4c",  x"4f",  x"53",  x"45",  x"cf", -- 1D88
         x"50",  x"45",  x"4e",  x"d2",  x"41",  x"4e",  x"44",  x"4f", -- 1D90
         x"4d",  x"49",  x"5a",  x"45",  x"d6",  x"47",  x"45",  x"54", -- 1D98
         x"24",  x"cc",  x"49",  x"4e",  x"45",  x"c3",  x"49",  x"52", -- 1DA0
         x"43",  x"4c",  x"45",  x"c3",  x"53",  x"52",  x"4c",  x"49", -- 1DA8
         x"4e",  x"80",  x"7d",  x"eb",  x"fd",  x"02",  x"06",  x"e7", -- 1DB0
         x"24",  x"ec",  x"65",  x"e7",  x"45",  x"e9",  x"6a",  x"e9", -- 1DB8
         x"9e",  x"e9",  x"b3",  x"e9",  x"89",  x"ea",  x"fa",  x"ea", -- 1DC0
         x"14",  x"eb",  x"48",  x"c3",  x"30",  x"eb",  x"98",  x"eb", -- 1DC8
         x"db",  x"eb",  x"0c",  x"ec",  x"3d",  x"ea",  x"48",  x"c3", -- 1DD0
         x"6c",  x"ea",  x"49",  x"eb",  x"a8",  x"ec",  x"99",  x"ec", -- 1DD8
         x"ac",  x"ec",  x"48",  x"c3",  x"f8",  x"ec",  x"39",  x"ed", -- 1DE0
         x"33",  x"ed",  x"48",  x"c3",  x"6e",  x"ed",  x"73",  x"ed", -- 1DE8
         x"00",  x"c0",  x"20",  x"8f",  x"00",  x"00",  x"00",  x"54", -- 1DF0
         x"80",  x"40",  x"20",  x"10",  x"08",  x"04",  x"02",  x"01", -- 1DF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"81",  x"ff", -- 1E00
         x"00",  x"00",  x"22",  x"72",  x"22",  x"3e",  x"00",  x"00", -- 1E08
         x"00",  x"00",  x"12",  x"32",  x"7e",  x"32",  x"12",  x"00", -- 1E10
         x"7e",  x"81",  x"b9",  x"a5",  x"b9",  x"a5",  x"b9",  x"81", -- 1E18
         x"55",  x"ff",  x"55",  x"ff",  x"55",  x"ff",  x"55",  x"ff", -- 1E20
         x"aa",  x"aa",  x"aa",  x"aa",  x"aa",  x"aa",  x"aa",  x"aa", -- 1E28
         x"ff",  x"00",  x"ff",  x"00",  x"ff",  x"00",  x"ff",  x"00", -- 1E30
         x"00",  x"00",  x"3c",  x"42",  x"42",  x"7e",  x"00",  x"00", -- 1E38
         x"00",  x"10",  x"30",  x"7e",  x"30",  x"10",  x"00",  x"00", -- 1E40
         x"00",  x"08",  x"0c",  x"7e",  x"0c",  x"08",  x"00",  x"00", -- 1E48
         x"00",  x"10",  x"10",  x"10",  x"7c",  x"38",  x"10",  x"00", -- 1E50
         x"08",  x"1c",  x"3e",  x"08",  x"08",  x"08",  x"08",  x"00", -- 1E58
         x"38",  x"30",  x"28",  x"08",  x"08",  x"08",  x"3e",  x"00", -- 1E60
         x"00",  x"00",  x"12",  x"32",  x"7e",  x"30",  x"10",  x"00", -- 1E68
         x"aa",  x"55",  x"aa",  x"55",  x"aa",  x"55",  x"aa",  x"55", -- 1E70
         x"3e",  x"7c",  x"7c",  x"3e",  x"3e",  x"7c",  x"f8",  x"f8", -- 1E78
         x"38",  x"30",  x"28",  x"04",  x"04",  x"04",  x"04",  x"00", -- 1E80
         x"7f",  x"08",  x"1c",  x"2a",  x"08",  x"08",  x"08",  x"00", -- 1E88
         x"00",  x"08",  x"08",  x"08",  x"2a",  x"1c",  x"08",  x"7f", -- 1E90
         x"7e",  x"81",  x"9d",  x"a1",  x"b9",  x"85",  x"85",  x"b9", -- 1E98
         x"00",  x"3c",  x"42",  x"5a",  x"5a",  x"42",  x"3c",  x"00", -- 1EA0
         x"88",  x"44",  x"22",  x"11",  x"88",  x"44",  x"22",  x"11", -- 1EA8
         x"00",  x"7f",  x"22",  x"72",  x"27",  x"22",  x"7f",  x"00", -- 1EB0
         x"11",  x"22",  x"44",  x"88",  x"11",  x"22",  x"44",  x"88", -- 1EB8
         x"00",  x"01",  x"09",  x"0d",  x"7f",  x"0d",  x"09",  x"01", -- 1EC0
         x"00",  x"90",  x"b0",  x"fe",  x"b0",  x"90",  x"00",  x"00", -- 1EC8
         x"00",  x"08",  x"7c",  x"06",  x"7c",  x"08",  x"00",  x"00", -- 1ED0
         x"cc",  x"cc",  x"33",  x"33",  x"cc",  x"cc",  x"33",  x"33", -- 1ED8
         x"7e",  x"81",  x"a1",  x"a1",  x"a1",  x"a1",  x"bd",  x"81", -- 1EE0
         x"7e",  x"81",  x"b9",  x"a5",  x"b9",  x"a5",  x"a5",  x"81", -- 1EE8
         x"7e",  x"81",  x"99",  x"a1",  x"a1",  x"a1",  x"99",  x"81", -- 1EF0
         x"00",  x"10",  x"3e",  x"60",  x"3e",  x"10",  x"00",  x"00", -- 1EF8
         x"3c",  x"42",  x"99",  x"a1",  x"a1",  x"99",  x"42",  x"3c", -- 1F00
         x"00",  x"00",  x"78",  x"0c",  x"7c",  x"cc",  x"76",  x"00", -- 1F08
         x"e0",  x"60",  x"7c",  x"66",  x"66",  x"66",  x"dc",  x"00", -- 1F10
         x"00",  x"00",  x"78",  x"cc",  x"c0",  x"cc",  x"78",  x"00", -- 1F18
         x"1c",  x"0c",  x"7c",  x"cc",  x"cc",  x"cc",  x"76",  x"00", -- 1F20
         x"00",  x"00",  x"78",  x"cc",  x"fc",  x"c0",  x"78",  x"00", -- 1F28
         x"38",  x"6c",  x"60",  x"f0",  x"60",  x"60",  x"f0",  x"00", -- 1F30
         x"00",  x"00",  x"76",  x"cc",  x"cc",  x"7c",  x"0c",  x"f8", -- 1F38
         x"e0",  x"60",  x"6c",  x"76",  x"66",  x"66",  x"e6",  x"00", -- 1F40
         x"30",  x"00",  x"70",  x"30",  x"30",  x"30",  x"fc",  x"00", -- 1F48
         x"0c",  x"00",  x"1c",  x"0c",  x"0c",  x"cc",  x"cc",  x"78", -- 1F50
         x"e0",  x"60",  x"66",  x"6c",  x"78",  x"6c",  x"e6",  x"00", -- 1F58
         x"70",  x"30",  x"30",  x"30",  x"30",  x"30",  x"fc",  x"00", -- 1F60
         x"00",  x"00",  x"cc",  x"fe",  x"fe",  x"d6",  x"c6",  x"00", -- 1F68
         x"00",  x"00",  x"f8",  x"cc",  x"cc",  x"cc",  x"cc",  x"00", -- 1F70
         x"00",  x"00",  x"78",  x"cc",  x"cc",  x"cc",  x"78",  x"00", -- 1F78
         x"00",  x"00",  x"dc",  x"66",  x"66",  x"7c",  x"60",  x"f0", -- 1F80
         x"00",  x"00",  x"76",  x"cc",  x"cc",  x"7c",  x"0c",  x"1e", -- 1F88
         x"00",  x"00",  x"dc",  x"76",  x"66",  x"60",  x"f0",  x"00", -- 1F90
         x"00",  x"00",  x"7c",  x"c0",  x"78",  x"0c",  x"f8",  x"00", -- 1F98
         x"10",  x"30",  x"7c",  x"30",  x"30",  x"34",  x"18",  x"00", -- 1FA0
         x"00",  x"00",  x"cc",  x"cc",  x"cc",  x"cc",  x"76",  x"00", -- 1FA8
         x"00",  x"00",  x"cc",  x"cc",  x"cc",  x"78",  x"30",  x"00", -- 1FB0
         x"00",  x"00",  x"c6",  x"d6",  x"fe",  x"fe",  x"6c",  x"00", -- 1FB8
         x"00",  x"00",  x"c6",  x"6c",  x"38",  x"6c",  x"c6",  x"00", -- 1FC0
         x"00",  x"00",  x"cc",  x"cc",  x"cc",  x"7c",  x"0c",  x"f8", -- 1FC8
         x"00",  x"00",  x"fc",  x"98",  x"30",  x"64",  x"fc",  x"00", -- 1FD0
         x"6c",  x"00",  x"78",  x"0c",  x"7c",  x"cc",  x"76",  x"00", -- 1FD8
         x"cc",  x"00",  x"78",  x"cc",  x"cc",  x"cc",  x"78",  x"00", -- 1FE0
         x"cc",  x"00",  x"cc",  x"cc",  x"cc",  x"cc",  x"76",  x"00", -- 1FE8
         x"3c",  x"66",  x"66",  x"6c",  x"66",  x"66",  x"6c",  x"f0", -- 1FF0
         x"ff",  x"81",  x"81",  x"81",  x"81",  x"81",  x"81",  x"ff"  -- 1FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
