library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_m012 is
    generic(
        ADDR_WIDTH   : integer := 13
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom_m012;

architecture rtl of rom_m012 is
    type rom8192x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom8192x8 := (
         x"00",  x"00",  x"3c",  x"66",  x"66",  x"66",  x"3b",  x"00", -- 0000
         x"00",  x"60",  x"60",  x"78",  x"6c",  x"6c",  x"78",  x"00", -- 0008
         x"00",  x"00",  x"3c",  x"66",  x"60",  x"66",  x"3c",  x"00", -- 0010
         x"00",  x"06",  x"06",  x"1e",  x"36",  x"36",  x"1e",  x"00", -- 0018
         x"00",  x"00",  x"38",  x"6c",  x"7c",  x"60",  x"38",  x"00", -- 0020
         x"00",  x"1e",  x"18",  x"7e",  x"18",  x"18",  x"18",  x"00", -- 0028
         x"00",  x"00",  x"3c",  x"66",  x"66",  x"3f",  x"06",  x"3c", -- 0030
         x"00",  x"60",  x"60",  x"6c",  x"76",  x"66",  x"66",  x"00", -- 0038
         x"00",  x"18",  x"00",  x"18",  x"18",  x"18",  x"18",  x"00", -- 0040
         x"00",  x"18",  x"00",  x"38",  x"18",  x"18",  x"18",  x"30", -- 0048
         x"00",  x"60",  x"66",  x"6c",  x"78",  x"6c",  x"66",  x"00", -- 0050
         x"00",  x"30",  x"30",  x"30",  x"30",  x"30",  x"18",  x"00", -- 0058
         x"00",  x"00",  x"36",  x"7f",  x"6b",  x"63",  x"63",  x"00", -- 0060
         x"00",  x"00",  x"7c",  x"66",  x"66",  x"66",  x"66",  x"00", -- 0068
         x"00",  x"00",  x"3c",  x"66",  x"66",  x"66",  x"3c",  x"00", -- 0070
         x"00",  x"00",  x"7c",  x"66",  x"66",  x"7c",  x"60",  x"60", -- 0078
         x"00",  x"00",  x"3c",  x"66",  x"66",  x"3e",  x"06",  x"06", -- 0080
         x"00",  x"00",  x"36",  x"38",  x"30",  x"30",  x"30",  x"00", -- 0088
         x"00",  x"00",  x"1c",  x"30",  x"1c",  x"06",  x"3c",  x"00", -- 0090
         x"00",  x"18",  x"18",  x"3c",  x"18",  x"18",  x"0c",  x"00", -- 0098
         x"00",  x"00",  x"66",  x"66",  x"66",  x"66",  x"3c",  x"00", -- 00A0
         x"00",  x"00",  x"66",  x"66",  x"3c",  x"3c",  x"18",  x"00", -- 00A8
         x"00",  x"00",  x"63",  x"63",  x"6b",  x"7f",  x"36",  x"00", -- 00B0
         x"00",  x"00",  x"66",  x"3c",  x"18",  x"3c",  x"66",  x"00", -- 00B8
         x"00",  x"00",  x"66",  x"3c",  x"18",  x"30",  x"60",  x"00", -- 00C0
         x"00",  x"00",  x"7e",  x"0c",  x"18",  x"30",  x"7e",  x"00", -- 00C8
         x"66",  x"00",  x"3c",  x"66",  x"66",  x"66",  x"3b",  x"00", -- 00D0
         x"66",  x"00",  x"3c",  x"64",  x"66",  x"66",  x"3c",  x"00", -- 00D8
         x"66",  x"00",  x"66",  x"66",  x"66",  x"66",  x"3c",  x"00", -- 00E0
         x"00",  x"1c",  x"34",  x"3c",  x"34",  x"3c",  x"30",  x"30", -- 00E8
         x"80",  x"40",  x"20",  x"10",  x"08",  x"04",  x"02",  x"01", -- 00F0
         x"3e",  x"00",  x"08",  x"08",  x"08",  x"2a",  x"1c",  x"08", -- 00F8
         x"c3",  x"3c",  x"66",  x"66",  x"7e",  x"66",  x"66",  x"00", -- 0100
         x"c3",  x"3c",  x"66",  x"66",  x"66",  x"66",  x"3c",  x"00", -- 0108
         x"81",  x"66",  x"66",  x"66",  x"66",  x"66",  x"3c",  x"00", -- 0110
         x"00",  x"7e",  x"42",  x"42",  x"42",  x"42",  x"7e",  x"00", -- 0118
         x"00",  x"18",  x"24",  x"42",  x"42",  x"24",  x"18",  x"00", -- 0120
         x"00",  x"18",  x"18",  x"24",  x"24",  x"42",  x"7e",  x"00", -- 0128
         x"00",  x"00",  x"00",  x"30",  x"49",  x"06",  x"00",  x"00", -- 0130
         x"a5",  x"eb",  x"c7",  x"d8",  x"d1",  x"da",  x"c1",  x"cf", -- 0138
         x"c0",  x"dc",  x"88",  x"e0",  x"86",  x"fe",  x"29",  x"c4", -- 0140
         x"d2",  x"a5",  x"a8",  x"a5",  x"ea",  x"cd",  x"ce",  x"cd", -- 0148
         x"c0",  x"c4",  x"92",  x"a8",  x"a4",  x"a5",  x"e3",  x"c7", -- 0150
         x"d8",  x"ce",  x"88",  x"a8",  x"fc",  x"cd",  x"d0",  x"dc", -- 0158
         x"a5",  x"a5",  x"a8",  x"a5",  x"ec",  x"cd",  x"c4",  x"cd", -- 0160
         x"dc",  x"cd",  x"88",  x"de",  x"c7",  x"c6",  x"88",  x"f2", -- 0168
         x"cd",  x"c1",  x"c4",  x"cd",  x"92",  x"a5",  x"a8",  x"88", -- 0170
         x"ca",  x"c1",  x"db",  x"92",  x"a5",  x"a8",  x"a5",  x"85", -- 0178
         x"88",  x"c1",  x"cb",  x"c0",  x"88",  x"db",  x"c7",  x"da", -- 0180
         x"dc",  x"c1",  x"cd",  x"da",  x"cd",  x"88",  x"85",  x"a5", -- 0188
         x"a8",  x"a5",  x"cd",  x"cc",  x"c1",  x"dc",  x"c1",  x"cd", -- 0190
         x"da",  x"cd",  x"c6",  x"a8",  x"a5",  x"fb",  x"d8",  x"cd", -- 0198
         x"c1",  x"cb",  x"c0",  x"cd",  x"da",  x"88",  x"d2",  x"dd", -- 01A0
         x"88",  x"c3",  x"c4",  x"cd",  x"c1",  x"c6",  x"a5",  x"a8", -- 01A8
         x"a4",  x"a5",  x"f2",  x"cd",  x"c1",  x"cb",  x"c0",  x"cd", -- 01B0
         x"c6",  x"c3",  x"cd",  x"dc",  x"dc",  x"cd",  x"88",  x"80", -- 01B8
         x"f3",  x"95",  x"cc",  x"c7",  x"c6",  x"dc",  x"88",  x"cb", -- 01C0
         x"c9",  x"da",  x"cd",  x"81",  x"92",  x"a5",  x"a8",  x"a4", -- 01C8
         x"de",  x"c7",  x"c6",  x"88",  x"f2",  x"cd",  x"c1",  x"c4", -- 01D0
         x"cd",  x"92",  x"a5",  x"a8",  x"a5",  x"f2",  x"cd",  x"c1", -- 01D8
         x"c4",  x"cd",  x"c6",  x"87",  x"fb",  x"cd",  x"c1",  x"dc", -- 01E0
         x"cd",  x"92",  x"a5",  x"a8",  x"a5",  x"ec",  x"da",  x"dd", -- 01E8
         x"cb",  x"c3",  x"88",  x"e2",  x"87",  x"e6",  x"92",  x"a5", -- 01F0
         x"a8",  x"a4",  x"e6",  x"c9",  x"c5",  x"cd",  x"92",  x"a5", -- 01F8
         x"a8",  x"a4",  x"e3",  x"c7",  x"d8",  x"ce",  x"d2",  x"cd", -- 0200
         x"c1",  x"c4",  x"cd",  x"c6",  x"92",  x"a5",  x"a8",  x"a4", -- 0208
         x"c5",  x"c1",  x"dc",  x"88",  x"8f",  x"84",  x"8f",  x"95", -- 0210
         x"e9",  x"fb",  x"eb",  x"e1",  x"e1",  x"84",  x"88",  x"db", -- 0218
         x"c7",  x"c6",  x"db",  x"dc",  x"88",  x"e0",  x"ed",  x"f0", -- 0220
         x"85",  x"ff",  x"cd",  x"da",  x"dc",  x"a5",  x"c9",  x"c4", -- 0228
         x"dc",  x"cd",  x"db",  x"88",  x"f2",  x"cd",  x"c1",  x"cb", -- 0230
         x"c0",  x"cd",  x"c6",  x"88",  x"a5",  x"a8",  x"a5",  x"c6", -- 0238
         x"cd",  x"dd",  x"cd",  x"db",  x"88",  x"f2",  x"cd",  x"c1", -- 0240
         x"cb",  x"c0",  x"cd",  x"c6",  x"88",  x"a5",  x"a8",  x"a5", -- 0248
         x"c6",  x"cd",  x"dd",  x"cd",  x"88",  x"e3",  x"cd",  x"dc", -- 0250
         x"dc",  x"cd",  x"92",  x"a5",  x"a8",  x"a5",  x"ee",  x"c1", -- 0258
         x"c4",  x"cd",  x"88",  x"a8",  x"88",  x"ea",  x"d1",  x"dc", -- 0260
         x"cd",  x"88",  x"c4",  x"c9",  x"c6",  x"cf",  x"a5",  x"c6", -- 0268
         x"c7",  x"cb",  x"c0",  x"88",  x"a8",  x"88",  x"ea",  x"d1", -- 0270
         x"dc",  x"cd",  x"88",  x"ce",  x"da",  x"cd",  x"c1",  x"a5", -- 0278
         x"a8",  x"a5",  x"d2",  x"dd",  x"c5",  x"88",  x"e9",  x"ca", -- 0280
         x"db",  x"c9",  x"dc",  x"d2",  x"92",  x"a5",  x"a8",  x"a5", -- 0288
         x"f2",  x"cd",  x"c1",  x"c4",  x"cd",  x"c6",  x"c4",  x"28", -- 0290
         x"c6",  x"cf",  x"cd",  x"92",  x"a5",  x"a8",  x"88",  x"f2", -- 0298
         x"cd",  x"c1",  x"cb",  x"c0",  x"cd",  x"c6",  x"a5",  x"88", -- 02A0
         x"f2",  x"cd",  x"c1",  x"c4",  x"cd",  x"c6",  x"a5",  x"fc", -- 02A8
         x"cd",  x"d0",  x"dc",  x"88",  x"a8",  x"88",  x"f2",  x"cd", -- 02B0
         x"c1",  x"c4",  x"cd",  x"c6",  x"a5",  x"a5",  x"a8",  x"a5", -- 02B8
         x"df",  x"c1",  x"da",  x"c3",  x"c4",  x"c1",  x"cb",  x"c0", -- 02C0
         x"97",  x"a5",  x"a8",  x"a4",  x"a5",  x"a8",  x"e7",  x"fb", -- 02C8
         x"a8",  x"a4",  x"88",  x"88",  x"88",  x"88",  x"8b",  x"8b", -- 02D0
         x"8b",  x"8b",  x"88",  x"fc",  x"cd",  x"d0",  x"dc",  x"de", -- 02D8
         x"cd",  x"da",  x"c9",  x"da",  x"ca",  x"cd",  x"c1",  x"dc", -- 02E0
         x"dd",  x"c6",  x"cf",  x"88",  x"8b",  x"8b",  x"8b",  x"8b", -- 02E8
         x"a5",  x"a5",  x"88",  x"88",  x"fe",  x"ed",  x"ea",  x"88", -- 02F0
         x"e5",  x"c1",  x"c3",  x"da",  x"c7",  x"cd",  x"c4",  x"cd", -- 02F8
         x"c3",  x"dc",  x"da",  x"c7",  x"c6",  x"c1",  x"c3",  x"88", -- 0300
         x"e5",  x"2a",  x"c0",  x"c4",  x"c0",  x"c9",  x"dd",  x"db", -- 0308
         x"cd",  x"c6",  x"a5",  x"fe",  x"cd",  x"da",  x"db",  x"c1", -- 0310
         x"c7",  x"c6",  x"88",  x"9a",  x"86",  x"9b",  x"a5",  x"85", -- 0318
         x"85",  x"85",  x"85",  x"85",  x"85",  x"85",  x"85",  x"85", -- 0320
         x"85",  x"85",  x"85",  x"85",  x"85",  x"85",  x"85",  x"85", -- 0328
         x"85",  x"85",  x"85",  x"85",  x"85",  x"85",  x"85",  x"85", -- 0330
         x"85",  x"85",  x"85",  x"85",  x"85",  x"85",  x"85",  x"85", -- 0338
         x"85",  x"a5",  x"a5",  x"e1",  x"92",  x"e1",  x"e6",  x"e1", -- 0340
         x"fc",  x"88",  x"88",  x"ee",  x"92",  x"ee",  x"e1",  x"e4", -- 0348
         x"ed",  x"f0",  x"88",  x"88",  x"fb",  x"92",  x"fb",  x"e7", -- 0350
         x"fa",  x"ed",  x"ec",  x"88",  x"88",  x"fc",  x"92",  x"fc", -- 0358
         x"ed",  x"f0",  x"e7",  x"fa",  x"a5",  x"a5",  x"fb",  x"fc", -- 0360
         x"e7",  x"f8",  x"88",  x"e0",  x"eb",  x"85",  x"eb",  x"e9", -- 0368
         x"e7",  x"fb",  x"a5",  x"a5",  x"a8",  x"a4",  x"88",  x"88", -- 0370
         x"88",  x"88",  x"88",  x"82",  x"82",  x"82",  x"82",  x"82", -- 0378
         x"82",  x"82",  x"82",  x"88",  x"fc",  x"ed",  x"f0",  x"e7", -- 0380
         x"fa",  x"88",  x"82",  x"82",  x"82",  x"82",  x"82",  x"82", -- 0388
         x"82",  x"82",  x"a5",  x"a5",  x"88",  x"88",  x"ed",  x"c1", -- 0390
         x"c6",  x"cf",  x"c9",  x"ca",  x"cd",  x"c6",  x"88",  x"88", -- 0398
         x"88",  x"88",  x"88",  x"e9",  x"c6",  x"d2",  x"cd",  x"c1", -- 03A0
         x"cf",  x"cd",  x"c6",  x"88",  x"88",  x"88",  x"88",  x"e9", -- 03A8
         x"dd",  x"db",  x"cf",  x"c9",  x"ca",  x"cd",  x"c6",  x"a5", -- 03B0
         x"a5",  x"e6",  x"92",  x"e6",  x"cd",  x"dd",  x"cd",  x"88", -- 03B8
         x"ec",  x"c9",  x"dc",  x"cd",  x"c1",  x"88",  x"88",  x"88", -- 03C0
         x"e0",  x"92",  x"e5",  x"cd",  x"c6",  x"dd",  x"88",  x"88", -- 03C8
         x"88",  x"88",  x"fa",  x"92",  x"fa",  x"c9",  x"c6",  x"cc", -- 03D0
         x"dc",  x"cd",  x"db",  x"dc",  x"a5",  x"fc",  x"92",  x"ec", -- 03D8
         x"c9",  x"dc",  x"cd",  x"c1",  x"c9",  x"c6",  x"ce",  x"c9", -- 03E0
         x"c6",  x"cf",  x"88",  x"88",  x"ee",  x"92",  x"ec",  x"c9", -- 03E8
         x"dc",  x"cd",  x"c1",  x"85",  x"88",  x"88",  x"cd",  x"92", -- 03F0
         x"ee",  x"c4",  x"c9",  x"dc",  x"dc",  x"cd",  x"da",  x"db", -- 03F8
         x"c9",  x"dc",  x"d2",  x"a5",  x"ea",  x"92",  x"ec",  x"c9", -- 0400
         x"dc",  x"cd",  x"c1",  x"cd",  x"c6",  x"cc",  x"cd",  x"88", -- 0408
         x"88",  x"88",  x"88",  x"88",  x"88",  x"df",  x"cd",  x"da", -- 0410
         x"dc",  x"cd",  x"88",  x"88",  x"88",  x"ed",  x"92",  x"ea", -- 0418
         x"c4",  x"c7",  x"cb",  x"c3",  x"db",  x"c9",  x"dc",  x"d2", -- 0420
         x"a5",  x"ef",  x"92",  x"ef",  x"cd",  x"c0",  x"cd",  x"88", -- 0428
         x"e9",  x"ca",  x"db",  x"c9",  x"dc",  x"d2",  x"85",  x"e6", -- 0430
         x"da",  x"86",  x"a5",  x"a5",  x"ea",  x"fa",  x"e3",  x"92", -- 0438
         x"e0",  x"c9",  x"dd",  x"d8",  x"dc",  x"c5",  x"cd",  x"c6", -- 0440
         x"dd",  x"a5",  x"c6",  x"84",  x"dc",  x"84",  x"ca",  x"84", -- 0448
         x"cf",  x"84",  x"d2",  x"88",  x"c5",  x"c1",  x"dc",  x"88", -- 0450
         x"c3",  x"c4",  x"cd",  x"c1",  x"c6",  x"cd",  x"c5",  x"88", -- 0458
         x"ee",  x"cd",  x"c6",  x"db",  x"dc",  x"cd",  x"da",  x"a5", -- 0460
         x"a5",  x"2d",  x"e9",  x"92",  x"e5",  x"c9",  x"cb",  x"c0", -- 0468
         x"cd",  x"88",  x"e9",  x"ca",  x"db",  x"c9",  x"dc",  x"d2", -- 0470
         x"88",  x"88",  x"2d",  x"fe",  x"92",  x"e4",  x"29",  x"db", -- 0478
         x"cb",  x"c0",  x"cd",  x"88",  x"e9",  x"ca",  x"db",  x"c9", -- 0480
         x"dc",  x"d2",  x"a5",  x"2c",  x"92",  x"da",  x"cd",  x"cb", -- 0488
         x"c0",  x"dc",  x"db",  x"ca",  x"2a",  x"c6",  x"cc",  x"c1", -- 0490
         x"cf",  x"88",  x"88",  x"88",  x"ff",  x"92",  x"e4",  x"29", -- 0498
         x"db",  x"cb",  x"c0",  x"cd",  x"88",  x"f2",  x"cd",  x"c1", -- 04A0
         x"cb",  x"c0",  x"cd",  x"c6",  x"88",  x"88",  x"22",  x"84", -- 04A8
         x"2d",  x"a5",  x"23",  x"92",  x"f2",  x"cd",  x"c6",  x"dc", -- 04B0
         x"da",  x"c1",  x"cd",  x"da",  x"cd",  x"88",  x"88",  x"88", -- 04B8
         x"88",  x"88",  x"88",  x"e4",  x"92",  x"e4",  x"29",  x"db", -- 04C0
         x"cb",  x"c0",  x"cd",  x"88",  x"f2",  x"cd",  x"c1",  x"cb", -- 04C8
         x"c0",  x"cd",  x"c6",  x"24",  x"84",  x"22",  x"84",  x"2d", -- 04D0
         x"a5",  x"21",  x"92",  x"fc",  x"c9",  x"ca",  x"dd",  x"c4", -- 04D8
         x"c4",  x"c1",  x"cd",  x"da",  x"cd",  x"88",  x"88",  x"88", -- 04E0
         x"88",  x"88",  x"ec",  x"92",  x"e4",  x"29",  x"db",  x"cb", -- 04E8
         x"c0",  x"cd",  x"88",  x"88",  x"88",  x"88",  x"88",  x"88", -- 04F0
         x"88",  x"22",  x"fc",  x"cd",  x"d0",  x"dc",  x"2d",  x"a5", -- 04F8
         x"f2",  x"92",  x"fb",  x"dd",  x"cb",  x"c0",  x"cd",  x"88", -- 0500
         x"e3",  x"cd",  x"dc",  x"dc",  x"cd",  x"88",  x"88",  x"88", -- 0508
         x"88",  x"f8",  x"92",  x"ec",  x"da",  x"dd",  x"cb",  x"c3", -- 0510
         x"cd",  x"88",  x"88",  x"88",  x"88",  x"88",  x"88",  x"88", -- 0518
         x"22",  x"fc",  x"cd",  x"d0",  x"dc",  x"2d",  x"a5",  x"88", -- 0520
         x"88",  x"ce",  x"c7",  x"da",  x"dc",  x"db",  x"cd",  x"dc", -- 0528
         x"d2",  x"cd",  x"c6",  x"88",  x"88",  x"88",  x"88",  x"88", -- 0530
         x"e5",  x"92",  x"fe",  x"cd",  x"da",  x"c4",  x"c9",  x"cf", -- 0538
         x"cd",  x"da",  x"cd",  x"88",  x"22",  x"fc",  x"cd",  x"d0", -- 0540
         x"dc",  x"22",  x"85",  x"96",  x"2d",  x"a5",  x"88",  x"88", -- 0548
         x"c5",  x"c1",  x"dc",  x"88",  x"fb",  x"c0",  x"c1",  x"ce", -- 0550
         x"dc",  x"88",  x"eb",  x"e4",  x"fa",  x"88",  x"88",  x"eb", -- 0558
         x"92",  x"e3",  x"c7",  x"d8",  x"c1",  x"cd",  x"da",  x"cd", -- 0560
         x"88",  x"88",  x"88",  x"22",  x"fc",  x"cd",  x"d0",  x"dc", -- 0568
         x"22",  x"85",  x"96",  x"2d",  x"a5",  x"a5",  x"a8",  x"a4", -- 0570
         x"88",  x"88",  x"88",  x"88",  x"88",  x"82",  x"82",  x"82", -- 0578
         x"82",  x"82",  x"82",  x"82",  x"82",  x"88",  x"fb",  x"e7", -- 0580
         x"fa",  x"ed",  x"ec",  x"88",  x"82",  x"82",  x"82",  x"82", -- 0588
         x"82",  x"82",  x"82",  x"82",  x"a5",  x"a5",  x"88",  x"ed", -- 0590
         x"c1",  x"c6",  x"cf",  x"c9",  x"ca",  x"cd",  x"c6",  x"88", -- 0598
         x"88",  x"88",  x"ee",  x"dd",  x"c6",  x"c3",  x"dc",  x"c1", -- 05A0
         x"c7",  x"c6",  x"cd",  x"c6",  x"88",  x"88",  x"88",  x"88", -- 05A8
         x"88",  x"e9",  x"dd",  x"db",  x"cf",  x"c9",  x"ca",  x"cd", -- 05B0
         x"c6",  x"a5",  x"a5",  x"e3",  x"92",  x"e3",  x"c7",  x"d8", -- 05B8
         x"ce",  x"88",  x"88",  x"88",  x"88",  x"88",  x"88",  x"fb", -- 05C0
         x"92",  x"fb",  x"c7",  x"da",  x"dc",  x"c1",  x"cd",  x"da", -- 05C8
         x"cd",  x"88",  x"88",  x"88",  x"88",  x"88",  x"e9",  x"92", -- 05D0
         x"e9",  x"dd",  x"db",  x"cf",  x"c9",  x"ca",  x"cd",  x"a5", -- 05D8
         x"fc",  x"92",  x"fc",  x"cd",  x"d0",  x"dc",  x"88",  x"88", -- 05E0
         x"88",  x"88",  x"88",  x"88",  x"f2",  x"92",  x"f2",  x"cd", -- 05E8
         x"c1",  x"cb",  x"c0",  x"cd",  x"c6",  x"db",  x"dd",  x"cb", -- 05F0
         x"c0",  x"cd",  x"88",  x"e0",  x"92",  x"e5",  x"cd",  x"c6", -- 05F8
         x"dd",  x"a5",  x"f5",  x"92",  x"fe",  x"cd",  x"da",  x"ca", -- 0600
         x"c1",  x"c6",  x"cc",  x"cd",  x"88",  x"88",  x"fd",  x"92", -- 0608
         x"fb",  x"dd",  x"cb",  x"c0",  x"cd",  x"88",  x"c7",  x"c0", -- 0610
         x"c6",  x"cd",  x"88",  x"88",  x"88",  x"ee",  x"92",  x"ec", -- 0618
         x"c9",  x"dc",  x"cd",  x"c1",  x"85",  x"a5",  x"ea",  x"fa", -- 0620
         x"e3",  x"92",  x"ea",  x"cd",  x"cd",  x"c6",  x"cc",  x"cd", -- 0628
         x"88",  x"88",  x"88",  x"88",  x"f2",  x"cd",  x"c1",  x"cb", -- 0630
         x"c0",  x"cd",  x"c6",  x"c3",  x"cd",  x"dc",  x"dc",  x"cd", -- 0638
         x"88",  x"88",  x"88",  x"df",  x"cd",  x"da",  x"dc",  x"cd", -- 0640
         x"a5",  x"88",  x"88",  x"88",  x"88",  x"88",  x"88",  x"88", -- 0648
         x"88",  x"88",  x"88",  x"88",  x"88",  x"ed",  x"92",  x"ed", -- 0650
         x"cc",  x"c1",  x"dc",  x"c1",  x"cd",  x"da",  x"cd",  x"a5", -- 0658
         x"a5",  x"c9",  x"84",  x"dd",  x"84",  x"d2",  x"88",  x"c7", -- 0660
         x"c0",  x"c6",  x"cd",  x"88",  x"f2",  x"cd",  x"c1",  x"c4", -- 0668
         x"cd",  x"c6",  x"85",  x"e6",  x"da",  x"86",  x"a5",  x"ea", -- 0670
         x"fa",  x"e3",  x"88",  x"a1",  x"e0",  x"c9",  x"dd",  x"d8", -- 0678
         x"dc",  x"c5",  x"cd",  x"c6",  x"dd",  x"a5",  x"a5",  x"ed", -- 0680
         x"cc",  x"c1",  x"dc",  x"c5",  x"c7",  x"cc",  x"cd",  x"a5", -- 0688
         x"e1",  x"e6",  x"fb",  x"84",  x"88",  x"ec",  x"ed",  x"e4", -- 0690
         x"84",  x"eb",  x"e4",  x"fa",  x"88",  x"dd",  x"db",  x"df", -- 0698
         x"86",  x"a5",  x"ed",  x"e6",  x"fc",  x"ed",  x"fa",  x"92", -- 06A0
         x"20",  x"ca",  x"cd",  x"da",  x"c6",  x"cd",  x"c0",  x"c5", -- 06A8
         x"cd",  x"a5",  x"ea",  x"fa",  x"e3",  x"92",  x"ea",  x"cd", -- 06B0
         x"cd",  x"c6",  x"cc",  x"cd",  x"a5",  x"a5",  x"a8",  x"a4", -- 06B8
         x"82",  x"82",  x"82",  x"82",  x"82",  x"82",  x"82",  x"82", -- 06C0
         x"82",  x"88",  x"ee",  x"e1",  x"e4",  x"ed",  x"f0",  x"88", -- 06C8
         x"82",  x"82",  x"82",  x"82",  x"82",  x"82",  x"82",  x"82", -- 06D0
         x"82",  x"a5",  x"a5",  x"a5",  x"88",  x"ee",  x"c1",  x"c4", -- 06D8
         x"cd",  x"88",  x"88",  x"88",  x"2e",  x"c6",  x"cc",  x"cd", -- 06E0
         x"da",  x"c6",  x"88",  x"88",  x"88",  x"ed",  x"da",  x"db", -- 06E8
         x"cd",  x"dc",  x"d2",  x"cd",  x"c6",  x"a5",  x"a5",  x"ee", -- 06F0
         x"92",  x"ff",  x"cd",  x"da",  x"dc",  x"cd",  x"88",  x"fb", -- 06F8
         x"85",  x"96",  x"fb",  x"e7",  x"fa",  x"ed",  x"ec",  x"88", -- 0700
         x"e3",  x"92",  x"e3",  x"cd",  x"dc",  x"dc",  x"cd",  x"c6", -- 0708
         x"a5",  x"e4",  x"92",  x"e4",  x"c9",  x"cc",  x"cd",  x"c6", -- 0710
         x"88",  x"fc",  x"85",  x"96",  x"fc",  x"ed",  x"f0",  x"e7", -- 0718
         x"fa",  x"88",  x"f2",  x"92",  x"f2",  x"cd",  x"c1",  x"cb", -- 0720
         x"c0",  x"cd",  x"c6",  x"a5",  x"e9",  x"92",  x"e9",  x"c6", -- 0728
         x"ce",  x"2a",  x"cf",  x"cd",  x"c6",  x"a5",  x"fa",  x"92", -- 0730
         x"fa",  x"cd",  x"dc",  x"dc",  x"cd",  x"c6",  x"a5",  x"a5", -- 0738
         x"ea",  x"fa",  x"e3",  x"92",  x"e0",  x"c9",  x"dd",  x"d8", -- 0740
         x"dc",  x"c5",  x"cd",  x"c6",  x"dd",  x"a5",  x"a5",  x"a8", -- 0748
         x"7f",  x"7f",  x"54",  x"45",  x"58",  x"54",  x"01",  x"f5", -- 0750
         x"c5",  x"d5",  x"e5",  x"cd",  x"1c",  x"c8",  x"3e",  x"80", -- 0758
         x"21",  x"00",  x"b9",  x"06",  x"0d",  x"36",  x"00",  x"23", -- 0760
         x"77",  x"23",  x"3c",  x"10",  x"f8",  x"00",  x"00",  x"00", -- 0768
         x"21",  x"00",  x"02",  x"23",  x"cb",  x"7c",  x"20",  x"08", -- 0770
         x"7e",  x"2f",  x"77",  x"be",  x"2f",  x"77",  x"28",  x"f3", -- 0778
         x"11",  x"68",  x"01",  x"b7",  x"ed",  x"52",  x"00",  x"00", -- 0780
         x"00",  x"00",  x"00",  x"00",  x"00",  x"22",  x"20",  x"01", -- 0788
         x"00",  x"00",  x"00",  x"cd",  x"58",  x"c8",  x"cd",  x"98", -- 0790
         x"c8",  x"3e",  x"01",  x"32",  x"00",  x"01",  x"00",  x"00", -- 0798
         x"cd",  x"4a",  x"c8",  x"cd",  x"e6",  x"c7",  x"21",  x"a6", -- 07A0
         x"c7",  x"e5",  x"c3",  x"a8",  x"dd",  x"06",  x"07",  x"21", -- 07A8
         x"4b",  x"c1",  x"cd",  x"29",  x"c8",  x"32",  x"22",  x"01", -- 07B0
         x"e6",  x"df",  x"2a",  x"23",  x"01",  x"22",  x"25",  x"01", -- 07B8
         x"eb",  x"be",  x"23",  x"28",  x"09",  x"23",  x"23",  x"10", -- 07C0
         x"f8",  x"c3",  x"45",  x"dd",  x"19",  x"c9",  x"7e",  x"23", -- 07C8
         x"66",  x"6f",  x"e9",  x"e1",  x"cd",  x"58",  x"c8",  x"21", -- 07D0
         x"cb",  x"c2",  x"c3",  x"f0",  x"dc",  x"e1",  x"d1",  x"c1", -- 07D8
         x"f1",  x"cd",  x"03",  x"f0",  x"12",  x"c9",  x"21",  x"d1", -- 07E0
         x"c2",  x"18",  x"0d",  x"21",  x"bf",  x"c6",  x"18",  x"08", -- 07E8
         x"21",  x"77",  x"c5",  x"18",  x"03",  x"21",  x"75",  x"c3", -- 07F0
         x"e5",  x"cd",  x"58",  x"c8",  x"e1",  x"cd",  x"0b",  x"c8", -- 07F8
         x"21",  x"00",  x"01",  x"11",  x"28",  x"1f",  x"18",  x"56", -- 0800
         x"c3",  x"30",  x"de",  x"7e",  x"ee",  x"a8",  x"b7",  x"c8", -- 0808
         x"23",  x"cd",  x"6b",  x"c8",  x"fe",  x"0d",  x"20",  x"f3", -- 0810
         x"3e",  x"0a",  x"18",  x"f5",  x"21",  x"f8",  x"be",  x"22", -- 0818
         x"a8",  x"b7",  x"21",  x"d0",  x"c0",  x"22",  x"ac",  x"b7", -- 0820
         x"c9",  x"cd",  x"0b",  x"c8",  x"cd",  x"31",  x"c8",  x"18", -- 0828
         x"3a",  x"e5",  x"cd",  x"03",  x"f0",  x"04",  x"fe",  x"41", -- 0830
         x"38",  x"0e",  x"fe",  x"5b",  x"38",  x"08",  x"fe",  x"61", -- 0838
         x"38",  x"06",  x"fe",  x"7b",  x"30",  x"02",  x"ee",  x"20", -- 0840
         x"e1",  x"c9",  x"1e",  x"06",  x"2e",  x"00",  x"3e",  x"02", -- 0848
         x"32",  x"81",  x"b7",  x"cd",  x"03",  x"f0",  x"0f",  x"c9", -- 0850
         x"21",  x"00",  x"00",  x"11",  x"28",  x"20",  x"22",  x"9c", -- 0858
         x"b7",  x"ed",  x"53",  x"9e",  x"b7",  x"c9",  x"cd",  x"4a", -- 0860
         x"c8",  x"3e",  x"0c",  x"cd",  x"03",  x"f0",  x"00",  x"c9", -- 0868
         x"db",  x"88",  x"cb",  x"d7",  x"d3",  x"88",  x"c9",  x"db", -- 0870
         x"88",  x"cb",  x"97",  x"18",  x"f7",  x"cd",  x"03",  x"f0", -- 0878
         x"24",  x"c9",  x"21",  x"bf",  x"c2",  x"cd",  x"29",  x"c8", -- 0880
         x"fe",  x"4a",  x"c0",  x"f5",  x"3e",  x"0d",  x"cd",  x"7d", -- 0888
         x"c8",  x"3e",  x"0a",  x"cd",  x"7d",  x"c8",  x"f1",  x"c9", -- 0890
         x"cd",  x"8b",  x"c8",  x"cd",  x"03",  x"f0",  x"20",  x"c9", -- 0898
         x"49",  x"58",  x"d9",  x"46",  x"47",  x"cf",  x"53",  x"67", -- 08A0
         x"ca",  x"54",  x"e8",  x"d0",  x"43",  x"08",  x"c8",  x"13", -- 08A8
         x"d3",  x"c7",  x"07",  x"e5",  x"c7",  x"e5",  x"ed",  x"5b", -- 08B0
         x"a0",  x"b7",  x"cd",  x"03",  x"f0",  x"32",  x"eb",  x"e1", -- 08B8
         x"c9",  x"22",  x"33",  x"01",  x"23",  x"cd",  x"0b",  x"c9", -- 08C0
         x"eb",  x"af",  x"57",  x"5f",  x"ed",  x"b1",  x"20",  x"03", -- 08C8
         x"13",  x"18",  x"f9",  x"ed",  x"53",  x"37",  x"01",  x"c9", -- 08D0
         x"e5",  x"1e",  x"01",  x"2e",  x"07",  x"cd",  x"4e",  x"c8", -- 08D8
         x"e1",  x"c3",  x"0b",  x"c8",  x"e5",  x"21",  x"00",  x"00", -- 08E0
         x"39",  x"af",  x"ed",  x"67",  x"f5",  x"ed",  x"67",  x"f5", -- 08E8
         x"23",  x"ed",  x"67",  x"f5",  x"ed",  x"67",  x"f5",  x"21", -- 08F0
         x"00",  x"00",  x"06",  x"04",  x"5d",  x"54",  x"29",  x"29", -- 08F8
         x"19",  x"29",  x"d1",  x"5a",  x"16",  x"00",  x"19",  x"10", -- 0900
         x"f3",  x"d1",  x"c9",  x"11",  x"01",  x"02",  x"b7",  x"ed", -- 0908
         x"52",  x"44",  x"4d",  x"c9",  x"c5",  x"d5",  x"e5",  x"af", -- 0910
         x"57",  x"06",  x"10",  x"29",  x"8f",  x"27",  x"5f",  x"7a", -- 0918
         x"8f",  x"27",  x"57",  x"cb",  x"11",  x"7b",  x"10",  x"f3", -- 0920
         x"eb",  x"3a",  x"3c",  x"01",  x"b7",  x"28",  x"05",  x"79", -- 0928
         x"cd",  x"03",  x"f0",  x"1c",  x"cd",  x"03",  x"f0",  x"1a", -- 0930
         x"3e",  x"20",  x"cd",  x"7d",  x"c8",  x"e1",  x"d1",  x"c1", -- 0938
         x"c9",  x"cd",  x"03",  x"f0",  x"1a",  x"3e",  x"20",  x"c3", -- 0940
         x"7d",  x"c8",  x"c5",  x"d5",  x"cd",  x"0b",  x"c8",  x"cd", -- 0948
         x"03",  x"f0",  x"17",  x"cd",  x"03",  x"f0",  x"22",  x"2a", -- 0950
         x"82",  x"b7",  x"cd",  x"e4",  x"c8",  x"eb",  x"2a",  x"37", -- 0958
         x"01",  x"b7",  x"ed",  x"52",  x"eb",  x"d1",  x"c1",  x"d0", -- 0960
         x"2a",  x"37",  x"01",  x"c9",  x"21",  x"78",  x"c1",  x"cd", -- 0968
         x"4a",  x"c9",  x"d8",  x"23",  x"c9",  x"11",  x"00",  x"02", -- 0970
         x"e5",  x"1a",  x"b7",  x"13",  x"20",  x"fb",  x"7c",  x"b5", -- 0978
         x"2b",  x"20",  x"f6",  x"e1",  x"c9",  x"e5",  x"d5",  x"c5", -- 0980
         x"21",  x"dc",  x"c1",  x"cd",  x"4a",  x"c9",  x"23",  x"22", -- 0988
         x"23",  x"01",  x"22",  x"2d",  x"01",  x"21",  x"ec",  x"c1", -- 0990
         x"cd",  x"29",  x"c8",  x"fe",  x"4a",  x"cd",  x"69",  x"c8", -- 0998
         x"20",  x"0a",  x"21",  x"4f",  x"c8",  x"cd",  x"03",  x"f0", -- 09A0
         x"1e",  x"cd",  x"8b",  x"c8",  x"c1",  x"d1",  x"e1",  x"c9", -- 09A8
         x"c5",  x"b7",  x"ed",  x"42",  x"e5",  x"c1",  x"e1",  x"c9", -- 09B0
         x"c5",  x"e5",  x"06",  x"07",  x"7e",  x"21",  x"59",  x"ca", -- 09B8
         x"be",  x"23",  x"28",  x"06",  x"23",  x"10",  x"f9",  x"e1", -- 09C0
         x"c1",  x"c9",  x"7e",  x"e1",  x"77",  x"c1",  x"c9",  x"c5", -- 09C8
         x"e5",  x"06",  x"07",  x"7e",  x"21",  x"66",  x"ca",  x"be", -- 09D0
         x"2b",  x"28",  x"ef",  x"2b",  x"10",  x"f9",  x"18",  x"e7", -- 09D8
         x"c1",  x"e1",  x"cb",  x"7e",  x"c4",  x"cf",  x"c9",  x"23", -- 09E0
         x"0b",  x"78",  x"b1",  x"20",  x"f5",  x"c3",  x"70",  x"c8", -- 09E8
         x"e5",  x"cd",  x"03",  x"f0",  x"0c",  x"30",  x"0c",  x"cd", -- 09F0
         x"03",  x"f0",  x"0e",  x"fe",  x"03",  x"28",  x"16",  x"fe", -- 09F8
         x"43",  x"20",  x"f4",  x"2a",  x"2d",  x"01",  x"2b",  x"7c", -- 0A00
         x"b5",  x"20",  x"07",  x"cd",  x"31",  x"c8",  x"b7",  x"2a", -- 0A08
         x"23",  x"01",  x"22",  x"2d",  x"01",  x"e1",  x"c9",  x"21", -- 0A10
         x"00",  x"00",  x"22",  x"37",  x"01",  x"22",  x"35",  x"01", -- 0A18
         x"21",  x"00",  x"02",  x"36",  x"00",  x"23",  x"22",  x"33", -- 0A20
         x"01",  x"c9",  x"21",  x"b0",  x"c1",  x"cd",  x"0b",  x"c8", -- 0A28
         x"2a",  x"20",  x"01",  x"23",  x"54",  x"5d",  x"cd",  x"31", -- 0A30
         x"c8",  x"fe",  x"01",  x"20",  x"0d",  x"e5",  x"b7",  x"ed", -- 0A38
         x"52",  x"e1",  x"28",  x"f2",  x"2b",  x"cd",  x"6b",  x"c8", -- 0A40
         x"18",  x"ec",  x"fe",  x"0d",  x"28",  x"08",  x"fe",  x"20", -- 0A48
         x"38",  x"e4",  x"77",  x"23",  x"18",  x"ef",  x"af",  x"77", -- 0A50
         x"c9",  x"80",  x"e1",  x"81",  x"ef",  x"82",  x"f5",  x"83", -- 0A58
         x"f3",  x"86",  x"c1",  x"87",  x"cf",  x"88",  x"d5",  x"2a", -- 0A60
         x"20",  x"01",  x"cd",  x"0b",  x"c9",  x"62",  x"6b",  x"3e", -- 0A68
         x"ff",  x"ed",  x"b1",  x"28",  x"05",  x"cd",  x"17",  x"ca", -- 0A70
         x"18",  x"12",  x"4e",  x"23",  x"46",  x"ed",  x"43",  x"35", -- 0A78
         x"01",  x"78",  x"a1",  x"3c",  x"ca",  x"c9",  x"c7",  x"2b", -- 0A80
         x"2b",  x"cd",  x"c1",  x"c8",  x"21",  x"19",  x"00",  x"22", -- 0A88
         x"23",  x"01",  x"cd",  x"f0",  x"c7",  x"af",  x"32",  x"3c", -- 0A90
         x"01",  x"21",  x"99",  x"ca",  x"e5",  x"c3",  x"60",  x"dd", -- 0A98
         x"06",  x"0c",  x"c3",  x"af",  x"c7",  x"3e",  x"0c",  x"32", -- 0AA0
         x"3c",  x"01",  x"cd",  x"6b",  x"c8",  x"21",  x"5d",  x"c2", -- 0AA8
         x"cd",  x"0b",  x"c8",  x"2a",  x"33",  x"01",  x"e5",  x"01", -- 0AB0
         x"00",  x"02",  x"b7",  x"ed",  x"42",  x"cd",  x"14",  x"c9", -- 0AB8
         x"21",  x"64",  x"c2",  x"cd",  x"0b",  x"c8",  x"2a",  x"20", -- 0AC0
         x"01",  x"c1",  x"b7",  x"ed",  x"42",  x"cd",  x"14",  x"c9", -- 0AC8
         x"af",  x"32",  x"3c",  x"01",  x"21",  x"75",  x"c2",  x"c3", -- 0AD0
         x"0b",  x"c8",  x"03",  x"fb",  x"ca",  x"53",  x"39",  x"cc", -- 0AD8
         x"54",  x"26",  x"cb",  x"41",  x"ca",  x"cb",  x"4b",  x"0c", -- 0AE0
         x"cb",  x"55",  x"32",  x"ce",  x"45",  x"3a",  x"cd",  x"46", -- 0AE8
         x"99",  x"cb",  x"5a",  x"32",  x"ce",  x"44",  x"c5",  x"ce", -- 0AF0
         x"48",  x"f0",  x"c7",  x"2a",  x"33",  x"01",  x"36",  x"ff", -- 0AF8
         x"ed",  x"5b",  x"35",  x"01",  x"23",  x"73",  x"23",  x"72", -- 0B00
         x"e1",  x"c3",  x"40",  x"dd",  x"21",  x"54",  x"c1",  x"cd", -- 0B08
         x"d8",  x"c8",  x"cd",  x"82",  x"c8",  x"20",  x"0c",  x"cd", -- 0B10
         x"17",  x"ca",  x"cd",  x"2f",  x"cb",  x"2a",  x"37",  x"01", -- 0B18
         x"22",  x"35",  x"01",  x"c3",  x"4a",  x"c8",  x"c3",  x"98", -- 0B20
         x"dd",  x"cd",  x"d8",  x"c8",  x"2a",  x"33",  x"01",  x"cd", -- 0B28
         x"b5",  x"c8",  x"06",  x"20",  x"cd",  x"31",  x"c8",  x"fe", -- 0B30
         x"03",  x"28",  x"e8",  x"fe",  x"0d",  x"28",  x"25",  x"fe", -- 0B38
         x"08",  x"28",  x"4a",  x"fe",  x"09",  x"28",  x"0c",  x"fe", -- 0B40
         x"1a",  x"28",  x"43",  x"fe",  x"1f",  x"28",  x"3f",  x"fe", -- 0B48
         x"20",  x"38",  x"e1",  x"cd",  x"6b",  x"c8",  x"fe",  x"5d", -- 0B50
         x"28",  x"0a",  x"10",  x"d8",  x"3e",  x"5d",  x"cd",  x"6b", -- 0B58
         x"c8",  x"00",  x"00",  x"00",  x"1a",  x"77",  x"23",  x"e5", -- 0B60
         x"d5",  x"ed",  x"5b",  x"20",  x"01",  x"b7",  x"ed",  x"52", -- 0B68
         x"d1",  x"e1",  x"30",  x"1f",  x"fe",  x"5d",  x"28",  x"10", -- 0B70
         x"13",  x"b7",  x"20",  x"e8",  x"22",  x"33",  x"01",  x"e5", -- 0B78
         x"2a",  x"37",  x"01",  x"23",  x"22",  x"37",  x"01",  x"e1", -- 0B80
         x"cd",  x"8b",  x"c8",  x"18",  x"a2",  x"04",  x"cd",  x"6b", -- 0B88
         x"c8",  x"18",  x"a1",  x"21",  x"9c",  x"c1",  x"cd",  x"0b", -- 0B90
         x"c8",  x"cd",  x"a5",  x"ca",  x"21",  x"55",  x"c1",  x"cd", -- 0B98
         x"0b",  x"c8",  x"2a",  x"35",  x"01",  x"e5",  x"cd",  x"14", -- 0BA0
         x"c9",  x"21",  x"a8",  x"c2",  x"cd",  x"0b",  x"c8",  x"2a", -- 0BA8
         x"37",  x"01",  x"2b",  x"cd",  x"14",  x"c9",  x"21",  x"b6", -- 0BB0
         x"c2",  x"cd",  x"0b",  x"c8",  x"3e",  x"63",  x"32",  x"22", -- 0BB8
         x"01",  x"21",  x"00",  x"00",  x"c1",  x"11",  x"01",  x"02", -- 0BC0
         x"18",  x"1e",  x"21",  x"cf",  x"c1",  x"cd",  x"4a",  x"c9", -- 0BC8
         x"e5",  x"e5",  x"cd",  x"75",  x"c9",  x"cd",  x"6c",  x"c9", -- 0BD0
         x"c1",  x"b7",  x"ed",  x"42",  x"e5",  x"c1",  x"e1",  x"da", -- 0BD8
         x"80",  x"dd",  x"ca",  x"80",  x"dd",  x"cd",  x"85",  x"c9", -- 0BE0
         x"cd",  x"f7",  x"cb",  x"ca",  x"98",  x"c8",  x"0b",  x"78", -- 0BE8
         x"b1",  x"ca",  x"98",  x"c8",  x"23",  x"18",  x"f1",  x"cd", -- 0BF0
         x"f0",  x"c9",  x"ca",  x"8b",  x"c8",  x"3a",  x"22",  x"01", -- 0BF8
         x"cb",  x"6f",  x"20",  x"1c",  x"cd",  x"14",  x"c9",  x"1a", -- 0C00
         x"13",  x"b7",  x"28",  x"27",  x"cd",  x"7d",  x"c8",  x"fe", -- 0C08
         x"5d",  x"20",  x"f4",  x"cd",  x"8b",  x"c8",  x"e5",  x"21", -- 0C10
         x"ff",  x"ff",  x"cd",  x"41",  x"c9",  x"e1",  x"18",  x"e7", -- 0C18
         x"1a",  x"13",  x"b7",  x"28",  x"0e",  x"fe",  x"5d",  x"20", -- 0C20
         x"05",  x"cd",  x"8b",  x"c8",  x"18",  x"f2",  x"cd",  x"7d", -- 0C28
         x"c8",  x"18",  x"ed",  x"cd",  x"8b",  x"c8",  x"fe",  x"01", -- 0C30
         x"c9",  x"cd",  x"82",  x"c8",  x"c0",  x"21",  x"7e",  x"c1", -- 0C38
         x"cd",  x"0b",  x"c8",  x"cd",  x"77",  x"c8",  x"2a",  x"35", -- 0C40
         x"01",  x"cd",  x"75",  x"c9",  x"ed",  x"53",  x"31",  x"01", -- 0C48
         x"d5",  x"2a",  x"33",  x"01",  x"b7",  x"ed",  x"52",  x"e5", -- 0C50
         x"e5",  x"c1",  x"eb",  x"cb",  x"7e",  x"c4",  x"b8",  x"c9", -- 0C58
         x"23",  x"0b",  x"78",  x"b1",  x"20",  x"f5",  x"2a",  x"33", -- 0C60
         x"01",  x"22",  x"25",  x"01",  x"2b",  x"af",  x"2b",  x"be", -- 0C68
         x"20",  x"fc",  x"23",  x"22",  x"27",  x"01",  x"af",  x"e5", -- 0C70
         x"ed",  x"5b",  x"31",  x"01",  x"b7",  x"ed",  x"52",  x"e1", -- 0C78
         x"ca",  x"e0",  x"c9",  x"2b",  x"2b",  x"be",  x"20",  x"fc", -- 0C80
         x"23",  x"22",  x"29",  x"01",  x"2a",  x"27",  x"01",  x"ed", -- 0C88
         x"5b",  x"29",  x"01",  x"7e",  x"e6",  x"5f",  x"47",  x"1a", -- 0C90
         x"e6",  x"5f",  x"b8",  x"28",  x"0d",  x"30",  x"19",  x"2a", -- 0C98
         x"27",  x"01",  x"22",  x"25",  x"01",  x"2a",  x"29",  x"01", -- 0CA0
         x"18",  x"c9",  x"b7",  x"28",  x"04",  x"23",  x"13",  x"18", -- 0CA8
         x"e2",  x"1a",  x"b7",  x"28",  x"ea",  x"be",  x"28",  x"f5", -- 0CB0
         x"2a",  x"27",  x"01",  x"ed",  x"4b",  x"29",  x"01",  x"cd", -- 0CB8
         x"b0",  x"c9",  x"c5",  x"ed",  x"5b",  x"33",  x"01",  x"ed", -- 0CC0
         x"b0",  x"2a",  x"29",  x"01",  x"ed",  x"5b",  x"25",  x"01", -- 0CC8
         x"7e",  x"e6",  x"5f",  x"47",  x"1a",  x"e6",  x"5f",  x"b8", -- 0CD0
         x"28",  x"1a",  x"30",  x"26",  x"2a",  x"33",  x"01",  x"ed", -- 0CD8
         x"5b",  x"25",  x"01",  x"b7",  x"ed",  x"52",  x"28",  x"30", -- 0CE0
         x"e5",  x"c1",  x"af",  x"d5",  x"e1",  x"ed",  x"b1",  x"22", -- 0CE8
         x"25",  x"01",  x"18",  x"d5",  x"b7",  x"28",  x"04",  x"23", -- 0CF0
         x"13",  x"18",  x"d5",  x"1a",  x"b7",  x"28",  x"dd",  x"be", -- 0CF8
         x"28",  x"f5",  x"2a",  x"25",  x"01",  x"ed",  x"4b",  x"27", -- 0D00
         x"01",  x"cd",  x"b0",  x"c9",  x"ed",  x"5b",  x"29",  x"01", -- 0D08
         x"ed",  x"b0",  x"c1",  x"2a",  x"33",  x"01",  x"18",  x"10", -- 0D10
         x"2a",  x"33",  x"01",  x"c1",  x"09",  x"ed",  x"4b",  x"27", -- 0D18
         x"01",  x"cd",  x"b0",  x"c9",  x"ed",  x"5b",  x"29",  x"01", -- 0D20
         x"ed",  x"b0",  x"2a",  x"29",  x"01",  x"e5",  x"af",  x"be", -- 0D28
         x"23",  x"20",  x"fc",  x"22",  x"25",  x"01",  x"e1",  x"c3", -- 0D30
         x"73",  x"cc",  x"21",  x"91",  x"c1",  x"cd",  x"0b",  x"c8", -- 0D38
         x"1e",  x"03",  x"2e",  x"07",  x"cd",  x"4e",  x"c8",  x"cd", -- 0D40
         x"31",  x"c8",  x"fe",  x"03",  x"ca",  x"66",  x"c8",  x"cd", -- 0D48
         x"6b",  x"c8",  x"fe",  x"0d",  x"20",  x"f1",  x"3e",  x"13", -- 0D50
         x"cd",  x"6b",  x"c8",  x"cd",  x"b5",  x"c8",  x"cd",  x"03", -- 0D58
         x"f0",  x"18",  x"da",  x"80",  x"dd",  x"3a",  x"96",  x"b7", -- 0D60
         x"fe",  x"04",  x"c2",  x"80",  x"dd",  x"13",  x"2a",  x"97", -- 0D68
         x"b7",  x"7c",  x"a5",  x"3c",  x"20",  x"07",  x"3e",  x"0b", -- 0D70
         x"cd",  x"6b",  x"c8",  x"18",  x"d9",  x"d5",  x"d5",  x"cd", -- 0D78
         x"e4",  x"c8",  x"d1",  x"eb",  x"2a",  x"37",  x"01",  x"2b", -- 0D80
         x"b7",  x"ed",  x"52",  x"eb",  x"d1",  x"da",  x"80",  x"dd", -- 0D88
         x"d5",  x"cd",  x"75",  x"c9",  x"ed",  x"53",  x"25",  x"01", -- 0D90
         x"23",  x"cd",  x"75",  x"c9",  x"ed",  x"53",  x"27",  x"01", -- 0D98
         x"e1",  x"ed",  x"5b",  x"33",  x"01",  x"23",  x"af",  x"be", -- 0DA0
         x"ca",  x"80",  x"dd",  x"e5",  x"e5",  x"01",  x"21",  x"00", -- 0DA8
         x"09",  x"af",  x"be",  x"0b",  x"2b",  x"28",  x"fb",  x"e1", -- 0DB0
         x"03",  x"03",  x"af",  x"b8",  x"20",  x"fa",  x"b9",  x"28", -- 0DB8
         x"f8",  x"ed",  x"b0",  x"2b",  x"7e",  x"fe",  x"5d",  x"e1", -- 0DC0
         x"20",  x"06",  x"01",  x"28",  x"00",  x"09",  x"18",  x"db", -- 0DC8
         x"af",  x"12",  x"2a",  x"25",  x"01",  x"ed",  x"5b",  x"33", -- 0DD0
         x"01",  x"af",  x"be",  x"1a",  x"77",  x"23",  x"13",  x"28", -- 0DD8
         x"20",  x"b7",  x"20",  x"f5",  x"e5",  x"2a",  x"33",  x"01", -- 0DE0
         x"ed",  x"5b",  x"27",  x"01",  x"cd",  x"0e",  x"c9",  x"e1", -- 0DE8
         x"28",  x"09",  x"38",  x"07",  x"eb",  x"ed",  x"b0",  x"ed", -- 0DF0
         x"53",  x"33",  x"01",  x"cd",  x"8b",  x"c8",  x"c3",  x"47", -- 0DF8
         x"cd",  x"b7",  x"28",  x"f7",  x"01",  x"00",  x"00",  x"2a", -- 0E00
         x"33",  x"01",  x"1a",  x"77",  x"23",  x"13",  x"03",  x"b7", -- 0E08
         x"20",  x"f8",  x"22",  x"33",  x"01",  x"e5",  x"09",  x"d1", -- 0E10
         x"eb",  x"c5",  x"e5",  x"ed",  x"4b",  x"27",  x"01",  x"cd", -- 0E18
         x"b0",  x"c9",  x"e1",  x"03",  x"ed",  x"b8",  x"2a",  x"33", -- 0E20
         x"01",  x"ed",  x"5b",  x"27",  x"01",  x"c1",  x"ed",  x"b0", -- 0E28
         x"18",  x"c9",  x"cd",  x"2a",  x"ca",  x"cd",  x"85",  x"c9", -- 0E30
         x"cd",  x"8b",  x"c8",  x"21",  x"ff",  x"ff",  x"22",  x"2b", -- 0E38
         x"01",  x"2a",  x"33",  x"01",  x"cd",  x"0b",  x"c9",  x"ed", -- 0E40
         x"43",  x"29",  x"01",  x"eb",  x"cd",  x"77",  x"c8",  x"22", -- 0E48
         x"31",  x"01",  x"e5",  x"af",  x"ed",  x"4b",  x"29",  x"01", -- 0E50
         x"ed",  x"b1",  x"ed",  x"43",  x"29",  x"01",  x"22",  x"27", -- 0E58
         x"01",  x"d1",  x"cd",  x"0e",  x"c9",  x"d5",  x"2a",  x"2b", -- 0E60
         x"01",  x"23",  x"22",  x"2b",  x"01",  x"ed",  x"5b",  x"37", -- 0E68
         x"01",  x"b7",  x"ed",  x"52",  x"e1",  x"28",  x"48",  x"ed", -- 0E70
         x"5b",  x"20",  x"01",  x"13",  x"1a",  x"ed",  x"b1",  x"28", -- 0E78
         x"0c",  x"3a",  x"22",  x"01",  x"cb",  x"47",  x"20",  x"23", -- 0E80
         x"2a",  x"27",  x"01",  x"18",  x"c2",  x"e5",  x"13",  x"1a", -- 0E88
         x"b7",  x"28",  x"10",  x"fe",  x"5b",  x"20",  x"03",  x"23", -- 0E90
         x"18",  x"f4",  x"ae",  x"e6",  x"df",  x"23",  x"28",  x"ee", -- 0E98
         x"e1",  x"18",  x"d4",  x"e1",  x"3a",  x"22",  x"01",  x"cb", -- 0EA0
         x"47",  x"20",  x"dd",  x"ed",  x"5b",  x"31",  x"01",  x"2a", -- 0EA8
         x"2b",  x"01",  x"cd",  x"70",  x"c8",  x"cd",  x"f7",  x"cb", -- 0EB0
         x"28",  x"08",  x"2a",  x"27",  x"01",  x"18",  x"8d",  x"cd", -- 0EB8
         x"70",  x"c8",  x"c3",  x"98",  x"c8",  x"21",  x"63",  x"c1", -- 0EC0
         x"cd",  x"4a",  x"c9",  x"cd",  x"75",  x"c9",  x"d5",  x"cd", -- 0EC8
         x"6c",  x"c9",  x"eb",  x"2a",  x"37",  x"01",  x"b7",  x"ed", -- 0ED0
         x"52",  x"e1",  x"d8",  x"28",  x"1a",  x"eb",  x"d5",  x"cd", -- 0ED8
         x"75",  x"c9",  x"e1",  x"e5",  x"b7",  x"ed",  x"52",  x"e1", -- 0EE0
         x"d2",  x"80",  x"dd",  x"e5",  x"2a",  x"33",  x"01",  x"cd", -- 0EE8
         x"0e",  x"c9",  x"c3",  x"70",  x"dd",  x"b0",  x"eb",  x"c3", -- 0EF0
         x"c1",  x"c8",  x"7f",  x"7f",  x"64",  x"01",  x"e5",  x"cd", -- 0EF8
         x"1c",  x"c8",  x"21",  x"1f",  x"00",  x"22",  x"23",  x"01", -- 0F00
         x"22",  x"2d",  x"01",  x"3e",  x"11",  x"cd",  x"6b",  x"c8", -- 0F08
         x"e1",  x"ed",  x"5b",  x"20",  x"01",  x"cd",  x"03",  x"f0", -- 0F10
         x"1a",  x"06",  x"20",  x"7e",  x"fe",  x"20",  x"30",  x"04", -- 0F18
         x"3e",  x"23",  x"18",  x"06",  x"fe",  x"8d",  x"38",  x"02", -- 0F20
         x"3e",  x"25",  x"cd",  x"6b",  x"c8",  x"23",  x"10",  x"eb", -- 0F28
         x"cd",  x"8b",  x"c8",  x"e5",  x"b7",  x"ed",  x"52",  x"e1", -- 0F30
         x"30",  x"05",  x"cd",  x"f0",  x"c9",  x"20",  x"d6",  x"3e", -- 0F38
         x"12",  x"cd",  x"6b",  x"c8",  x"c3",  x"8b",  x"c8",  x"cd", -- 0F40
         x"eb",  x"c7",  x"21",  x"4a",  x"cf",  x"e5",  x"06",  x"0a", -- 0F48
         x"c3",  x"b8",  x"dd",  x"c3",  x"af",  x"c7",  x"48",  x"eb", -- 0F50
         x"c7",  x"4b",  x"1d",  x"d0",  x"41",  x"cb",  x"d0",  x"4c", -- 0F58
         x"c2",  x"d0",  x"52",  x"99",  x"cf",  x"53",  x"be",  x"cf", -- 0F60
         x"54",  x"cd",  x"cf",  x"5a",  x"00",  x"d0",  x"46",  x"83", -- 0F68
         x"cf",  x"03",  x"74",  x"cf",  x"e1",  x"c3",  x"a3",  x"c7", -- 0F70
         x"01",  x"ff",  x"ff",  x"3e",  x"ff",  x"21",  x"00",  x"02", -- 0F78
         x"ed",  x"b1",  x"c9",  x"cd",  x"a5",  x"ca",  x"cd",  x"78", -- 0F80
         x"cf",  x"7e",  x"23",  x"a6",  x"21",  x"b4",  x"d0",  x"fe", -- 0F88
         x"ff",  x"20",  x"03",  x"21",  x"bb",  x"d0",  x"c3",  x"0b", -- 0F90
         x"c8",  x"21",  x"f9",  x"c1",  x"cd",  x"0b",  x"c8",  x"cd", -- 0F98
         x"03",  x"f0",  x"17",  x"d5",  x"3e",  x"02",  x"32",  x"81", -- 0FA0
         x"b7",  x"21",  x"00",  x"02",  x"22",  x"82",  x"b7",  x"cd", -- 0FA8
         x"78",  x"cf",  x"23",  x"23",  x"23",  x"22",  x"84",  x"b7", -- 0FB0
         x"e1",  x"cd",  x"03",  x"f0",  x"36",  x"c9",  x"21",  x"01", -- 0FB8
         x"c2",  x"cd",  x"4a",  x"c9",  x"e5",  x"cd",  x"78",  x"cf", -- 0FC0
         x"d1",  x"73",  x"23",  x"72",  x"c9",  x"cd",  x"78",  x"cf", -- 0FC8
         x"36",  x"ff",  x"23",  x"36",  x"ff",  x"c9",  x"cd",  x"31", -- 0FD0
         x"c8",  x"c3",  x"6b",  x"c8",  x"cd",  x"0b",  x"c8",  x"cd", -- 0FD8
         x"d6",  x"cf",  x"fe",  x"2c",  x"20",  x"04",  x"cd",  x"d6", -- 0FE0
         x"cf",  x"c9",  x"11",  x"3b",  x"01",  x"12",  x"cd",  x"d6", -- 0FE8
         x"cf",  x"13",  x"12",  x"1b",  x"cd",  x"03",  x"f0",  x"18", -- 0FF0
         x"38",  x"04",  x"3a",  x"97",  x"b7",  x"c9",  x"e1",  x"c9", -- 0FF8
         x"21",  x"0f",  x"c2",  x"cd",  x"dc",  x"cf",  x"4f",  x"21", -- 1000
         x"3e",  x"c2",  x"cd",  x"dc",  x"cf",  x"47",  x"21",  x"00", -- 1008
         x"02",  x"23",  x"3e",  x"ff",  x"be",  x"c8",  x"79",  x"be", -- 1010
         x"20",  x"f7",  x"70",  x"18",  x"f4",  x"cd",  x"78",  x"cf", -- 1018
         x"23",  x"23",  x"23",  x"22",  x"33",  x"01",  x"cd",  x"2a", -- 1020
         x"ca",  x"21",  x"4f",  x"c2",  x"cd",  x"0b",  x"c8",  x"21", -- 1028
         x"3b",  x"01",  x"cd",  x"34",  x"ca",  x"21",  x"3b",  x"01", -- 1030
         x"af",  x"47",  x"04",  x"be",  x"23",  x"20",  x"fb",  x"2a", -- 1038
         x"20",  x"01",  x"23",  x"05",  x"be",  x"20",  x"fb",  x"21", -- 1040
         x"00",  x"02",  x"ed",  x"5b",  x"20",  x"01",  x"13",  x"1a", -- 1048
         x"be",  x"23",  x"28",  x"06",  x"3e",  x"ff",  x"be",  x"c8", -- 1050
         x"18",  x"f5",  x"e5",  x"13",  x"1a",  x"b7",  x"28",  x"0e", -- 1058
         x"fe",  x"5b",  x"20",  x"03",  x"23",  x"18",  x"f4",  x"be", -- 1060
         x"23",  x"28",  x"f0",  x"e1",  x"18",  x"dc",  x"e1",  x"2b", -- 1068
         x"78",  x"b7",  x"20",  x"0c",  x"11",  x"3b",  x"01",  x"1a", -- 1070
         x"b7",  x"28",  x"cf",  x"77",  x"23",  x"13",  x"18",  x"f7", -- 1078
         x"ed",  x"5b",  x"33",  x"01",  x"eb",  x"b7",  x"ed",  x"52", -- 1080
         x"eb",  x"fe",  x"7f",  x"c5",  x"e5",  x"48",  x"06",  x"00", -- 1088
         x"38",  x"12",  x"e5",  x"af",  x"91",  x"4f",  x"09",  x"42", -- 1090
         x"4b",  x"d1",  x"ed",  x"b0",  x"ed",  x"53",  x"33",  x"01", -- 1098
         x"e1",  x"c1",  x"18",  x"d0",  x"2a",  x"33",  x"01",  x"e5", -- 10A0
         x"09",  x"22",  x"33",  x"01",  x"42",  x"4b",  x"d1",  x"eb", -- 10A8
         x"ed",  x"b8",  x"18",  x"ec",  x"fb",  x"e7",  x"fa",  x"ed", -- 10B0
         x"ec",  x"a5",  x"a8",  x"fc",  x"ed",  x"f0",  x"e7",  x"fa", -- 10B8
         x"a5",  x"a8",  x"af",  x"32",  x"81",  x"b7",  x"cd",  x"03", -- 10C0
         x"f0",  x"10",  x"c9",  x"cd",  x"78",  x"cf",  x"2b",  x"11", -- 10C8
         x"00",  x"02",  x"b7",  x"ed",  x"52",  x"22",  x"82",  x"b7", -- 10D0
         x"3e",  x"01",  x"cd",  x"c3",  x"d0",  x"3e",  x"ff",  x"2a", -- 10D8
         x"20",  x"01",  x"77",  x"2b",  x"77",  x"2b",  x"77",  x"c9", -- 10E0
         x"cd",  x"58",  x"c8",  x"af",  x"32",  x"3c",  x"01",  x"2a", -- 10E8
         x"20",  x"01",  x"11",  x"02",  x"02",  x"cd",  x"0e",  x"c9", -- 10F0
         x"d5",  x"e1",  x"2b",  x"3e",  x"ff",  x"ed",  x"b1",  x"28", -- 10F8
         x"01",  x"eb",  x"2b",  x"22",  x"33",  x"01",  x"3e",  x"3c", -- 1100
         x"32",  x"35",  x"01",  x"21",  x"ff",  x"ff",  x"22",  x"37", -- 1108
         x"01",  x"cd",  x"f5",  x"c7",  x"c3",  x"c8",  x"dd",  x"cd", -- 1110
         x"29",  x"c8",  x"32",  x"22",  x"01",  x"e6",  x"df",  x"21", -- 1118
         x"14",  x"d1",  x"e5",  x"21",  x"11",  x"d8",  x"06",  x"0c", -- 1120
         x"be",  x"23",  x"28",  x"07",  x"23",  x"23",  x"10",  x"f8", -- 1128
         x"c3",  x"c9",  x"c7",  x"7e",  x"23",  x"66",  x"6f",  x"e5", -- 1130
         x"78",  x"fe",  x"01",  x"38",  x"11",  x"fe",  x"09",  x"38", -- 1138
         x"0f",  x"3a",  x"22",  x"01",  x"cb",  x"6f",  x"cd",  x"69", -- 1140
         x"d1",  x"1e",  x"00",  x"c3",  x"30",  x"dd",  x"e1",  x"e9", -- 1148
         x"fe",  x"03",  x"cd",  x"69",  x"d1",  x"cd",  x"5f",  x"d1", -- 1150
         x"18",  x"f4",  x"2e",  x"06",  x"c3",  x"4e",  x"c8",  x"1e", -- 1158
         x"07",  x"2e",  x"00",  x"cd",  x"4e",  x"c8",  x"c3",  x"69", -- 1160
         x"c8",  x"20",  x"07",  x"3e",  x"1f",  x"21",  x"b0",  x"04", -- 1168
         x"18",  x"05",  x"3e",  x"07",  x"21",  x"f0",  x"00",  x"32", -- 1170
         x"9f",  x"b7",  x"22",  x"39",  x"01",  x"c9",  x"cd",  x"a5", -- 1178
         x"ca",  x"21",  x"90",  x"c2",  x"cd",  x"0b",  x"c8",  x"3a", -- 1180
         x"35",  x"01",  x"26",  x"00",  x"6f",  x"cd",  x"14",  x"c9", -- 1188
         x"21",  x"45",  x"c2",  x"c3",  x"2f",  x"df",  x"cd",  x"a0", -- 1190
         x"d4",  x"21",  x"ff",  x"ff",  x"22",  x"35",  x"01",  x"c3", -- 1198
         x"fb",  x"ca",  x"21",  x"81",  x"c2",  x"cd",  x"4a",  x"c9", -- 11A0
         x"e5",  x"c1",  x"21",  x"00",  x"02",  x"af",  x"23",  x"be", -- 11A8
         x"20",  x"fc",  x"e5",  x"ed",  x"5b",  x"33",  x"01",  x"1b", -- 11B0
         x"b7",  x"ed",  x"52",  x"e1",  x"30",  x"07",  x"0b",  x"78", -- 11B8
         x"b1",  x"20",  x"ea",  x"18",  x"0c",  x"2a",  x"33",  x"01", -- 11C0
         x"c3",  x"ca",  x"d2",  x"cd",  x"da",  x"d4",  x"21",  x"00", -- 11C8
         x"02",  x"e5",  x"2a",  x"a4",  x"b7",  x"22",  x"1e",  x"01", -- 11D0
         x"21",  x"40",  x"d8",  x"22",  x"a4",  x"b7",  x"cd",  x"4b", -- 11D8
         x"d8",  x"cd",  x"69",  x"c8",  x"cd",  x"4f",  x"d8",  x"e1", -- 11E0
         x"ed",  x"5b",  x"33",  x"01",  x"23",  x"22",  x"31",  x"01", -- 11E8
         x"18",  x"05",  x"7e",  x"cd",  x"6b",  x"c8",  x"23",  x"e5", -- 11F0
         x"b7",  x"ed",  x"52",  x"e1",  x"28",  x"23",  x"b7",  x"cc", -- 11F8
         x"8b",  x"c8",  x"cd",  x"26",  x"d2",  x"20",  x"eb",  x"eb", -- 1200
         x"e5",  x"cd",  x"0e",  x"c9",  x"e1",  x"ed",  x"5b",  x"20", -- 1208
         x"01",  x"1b",  x"2b",  x"ed",  x"b8",  x"13",  x"ed",  x"53", -- 1210
         x"2f",  x"01",  x"3e",  x"10",  x"cd",  x"6b",  x"c8",  x"18", -- 1218
         x"0f",  x"cd",  x"e9",  x"d4",  x"18",  x"f4",  x"3a",  x"a1", -- 1220
         x"b7",  x"3c",  x"47",  x"3a",  x"9f",  x"b7",  x"90",  x"c9", -- 1228
         x"c3",  x"90",  x"de",  x"fe",  x"03",  x"28",  x"38",  x"fe", -- 1230
         x"0c",  x"28",  x"34",  x"fe",  x"13",  x"28",  x"30",  x"fe", -- 1238
         x"11",  x"ca",  x"c7",  x"d2",  x"fe",  x"12",  x"ca",  x"d8", -- 1240
         x"d2",  x"fe",  x"0b",  x"28",  x"5d",  x"fe",  x"1a",  x"28", -- 1248
         x"2a",  x"fe",  x"0d",  x"28",  x"15",  x"fe",  x"0f",  x"ca", -- 1250
         x"8c",  x"d4",  x"fe",  x"85",  x"ca",  x"f3",  x"d2",  x"cd", -- 1258
         x"6b",  x"c8",  x"cd",  x"26",  x"d2",  x"cc",  x"14",  x"d5", -- 1260
         x"18",  x"c6",  x"cd",  x"8b",  x"c8",  x"18",  x"f3",  x"cd", -- 1268
         x"f6",  x"d4",  x"2a",  x"1e",  x"01",  x"22",  x"a4",  x"b7", -- 1270
         x"c3",  x"5f",  x"d1",  x"cd",  x"6b",  x"c8",  x"2a",  x"a0", -- 1278
         x"b7",  x"e5",  x"3a",  x"9f",  x"b7",  x"3d",  x"57",  x"1e", -- 1280
         x"00",  x"cd",  x"03",  x"f0",  x"32",  x"7e",  x"b7",  x"28", -- 1288
         x"13",  x"ed",  x"53",  x"a0",  x"b7",  x"2a",  x"2f",  x"01", -- 1290
         x"77",  x"2b",  x"36",  x"00",  x"22",  x"2f",  x"01",  x"3e", -- 1298
         x"02",  x"cd",  x"6b",  x"c8",  x"e1",  x"22",  x"a0",  x"b7", -- 12A0
         x"18",  x"86",  x"3a",  x"a1",  x"b7",  x"b7",  x"3e",  x"0b", -- 12A8
         x"c2",  x"5f",  x"d2",  x"cd",  x"e0",  x"d2",  x"cd",  x"e9", -- 12B0
         x"d2",  x"e5",  x"11",  x"00",  x"02",  x"b7",  x"ed",  x"52", -- 12B8
         x"e1",  x"da",  x"ce",  x"d1",  x"c3",  x"d1",  x"d1",  x"cd", -- 12C0
         x"e0",  x"d2",  x"3a",  x"9f",  x"b7",  x"3d",  x"47",  x"c5", -- 12C8
         x"cd",  x"e9",  x"d2",  x"c1",  x"10",  x"f9",  x"18",  x"e1", -- 12D0
         x"cd",  x"f6",  x"d4",  x"2a",  x"31",  x"01",  x"18",  x"d6", -- 12D8
         x"2a",  x"31",  x"01",  x"e5",  x"cd",  x"f6",  x"d4",  x"e1", -- 12E0
         x"c9",  x"01",  x"27",  x"00",  x"2b",  x"2b",  x"af",  x"ed", -- 12E8
         x"b9",  x"23",  x"c9",  x"cd",  x"6b",  x"c8",  x"cd",  x"f6", -- 12F0
         x"d4",  x"cd",  x"31",  x"c8",  x"b7",  x"28",  x"fa",  x"cb", -- 12F8
         x"af",  x"32",  x"2b",  x"01",  x"fe",  x"44",  x"ca",  x"c4", -- 1300
         x"d3",  x"fe",  x"50",  x"ca",  x"68",  x"d5",  x"fe",  x"43", -- 1308
         x"28",  x"30",  x"fe",  x"4d",  x"28",  x"2c",  x"fe",  x"41", -- 1310
         x"28",  x"0f",  x"fe",  x"56",  x"28",  x"12",  x"cd",  x"5f", -- 1318
         x"d1",  x"c3",  x"80",  x"dd",  x"2a",  x"29",  x"01",  x"18", -- 1320
         x"8d",  x"cd",  x"d0",  x"d4",  x"af",  x"77",  x"18",  x"86", -- 1328
         x"cd",  x"d0",  x"d4",  x"e5",  x"23",  x"23",  x"e5",  x"22", -- 1330
         x"29",  x"01",  x"eb",  x"cd",  x"f0",  x"d4",  x"e1",  x"d1", -- 1338
         x"18",  x"5f",  x"cd",  x"e4",  x"d3",  x"28",  x"d7",  x"2a", -- 1340
         x"27",  x"01",  x"ed",  x"5b",  x"25",  x"01",  x"cd",  x"0e", -- 1348
         x"c9",  x"0b",  x"78",  x"b1",  x"28",  x"c8",  x"2a",  x"33", -- 1350
         x"01",  x"e5",  x"09",  x"e5",  x"ed",  x"5b",  x"20",  x"01", -- 1358
         x"b7",  x"ed",  x"52",  x"d1",  x"e1",  x"30",  x"46",  x"3a", -- 1360
         x"2c",  x"01",  x"fe",  x"8a",  x"cc",  x"b3",  x"d3",  x"ed", -- 1368
         x"53",  x"33",  x"01",  x"c5",  x"e5",  x"ed",  x"4b",  x"29", -- 1370
         x"01",  x"b7",  x"ed",  x"42",  x"e5",  x"c1",  x"e1",  x"03", -- 1378
         x"ed",  x"b8",  x"c1",  x"c5",  x"ed",  x"5b",  x"29",  x"01", -- 1380
         x"2a",  x"25",  x"01",  x"23",  x"ed",  x"b0",  x"c1",  x"3a", -- 1388
         x"2b",  x"01",  x"fe",  x"43",  x"28",  x"11",  x"ed",  x"5b", -- 1390
         x"27",  x"01",  x"cd",  x"f0",  x"d4",  x"2a",  x"25",  x"01", -- 1398
         x"eb",  x"ed",  x"b0",  x"ed",  x"53",  x"33",  x"01",  x"cd", -- 13A0
         x"a5",  x"d4",  x"c3",  x"24",  x"d3",  x"cd",  x"5f",  x"d1", -- 13A8
         x"c3",  x"4d",  x"d5",  x"e5",  x"2a",  x"25",  x"01",  x"09", -- 13B0
         x"22",  x"25",  x"01",  x"2a",  x"27",  x"01",  x"09",  x"22", -- 13B8
         x"27",  x"01",  x"e1",  x"c9",  x"cd",  x"e3",  x"d3",  x"ca", -- 13C0
         x"1e",  x"d3",  x"ed",  x"5b",  x"29",  x"01",  x"13",  x"cd", -- 13C8
         x"f0",  x"d4",  x"2a",  x"27",  x"01",  x"eb",  x"ed",  x"b0", -- 13D0
         x"1b",  x"ed",  x"53",  x"33",  x"01",  x"2a",  x"27",  x"01", -- 13D8
         x"c3",  x"b6",  x"d2",  x"af",  x"11",  x"00",  x"02",  x"cd", -- 13E0
         x"f0",  x"d4",  x"eb",  x"23",  x"b7",  x"28",  x"3a",  x"7e", -- 13E8
         x"fe",  x"8a",  x"28",  x"2d",  x"fe",  x"85",  x"28",  x"07", -- 13F0
         x"23",  x"0b",  x"78",  x"b1",  x"c8",  x"18",  x"f0",  x"22", -- 13F8
         x"29",  x"01",  x"23",  x"0b",  x"78",  x"b1",  x"c8",  x"7e", -- 1400
         x"fe",  x"8a",  x"20",  x"f6",  x"22",  x"25",  x"01",  x"23", -- 1408
         x"0b",  x"78",  x"b1",  x"c8",  x"7e",  x"fe",  x"8a",  x"20", -- 1410
         x"f6",  x"22",  x"27",  x"01",  x"32",  x"2c",  x"01",  x"b7", -- 1418
         x"c9",  x"22",  x"25",  x"01",  x"23",  x"0b",  x"78",  x"b1", -- 1420
         x"c8",  x"7e",  x"fe",  x"8a",  x"20",  x"f6",  x"22",  x"27", -- 1428
         x"01",  x"23",  x"0b",  x"78",  x"b1",  x"c8",  x"7e",  x"fe", -- 1430
         x"85",  x"20",  x"f6",  x"22",  x"29",  x"01",  x"18",  x"dc", -- 1438
         x"cd",  x"2a",  x"ca",  x"01",  x"00",  x"02",  x"3e",  x"ff", -- 1440
         x"32",  x"25",  x"01",  x"2a",  x"33",  x"01",  x"c5",  x"b7", -- 1448
         x"ed",  x"42",  x"e5",  x"c1",  x"e1",  x"ed",  x"5b",  x"20", -- 1450
         x"01",  x"13",  x"04",  x"c5",  x"41",  x"23",  x"1a",  x"ae", -- 1458
         x"e6",  x"df",  x"28",  x"0a",  x"10",  x"f7",  x"c1",  x"0e", -- 1460
         x"00",  x"10",  x"f0",  x"c3",  x"5f",  x"d1",  x"d5",  x"e5", -- 1468
         x"c5",  x"13",  x"23",  x"1a",  x"b7",  x"28",  x"0e",  x"fe", -- 1470
         x"5b",  x"28",  x"f6",  x"ae",  x"e6",  x"df",  x"28",  x"f1", -- 1478
         x"c1",  x"e1",  x"d1",  x"18",  x"df",  x"c1",  x"e1",  x"d1", -- 1480
         x"c1",  x"c3",  x"b6",  x"d2",  x"cd",  x"f6",  x"d4",  x"3a", -- 1488
         x"25",  x"01",  x"3c",  x"c2",  x"5f",  x"d1",  x"2a",  x"31", -- 1490
         x"01",  x"cd",  x"e9",  x"d2",  x"e5",  x"c1",  x"18",  x"a6", -- 1498
         x"3e",  x"8c",  x"cd",  x"ac",  x"d4",  x"3e",  x"85",  x"cd", -- 14A0
         x"ac",  x"d4",  x"3e",  x"8a",  x"11",  x"01",  x"02",  x"cd", -- 14A8
         x"f0",  x"d4",  x"eb",  x"ed",  x"b1",  x"c0",  x"eb",  x"cd", -- 14B0
         x"f0",  x"d4",  x"d5",  x"e1",  x"1b",  x"d5",  x"ed",  x"b0", -- 14B8
         x"ed",  x"53",  x"33",  x"01",  x"d1",  x"18",  x"e8",  x"cd", -- 14C0
         x"03",  x"f0",  x"1a",  x"3e",  x"20",  x"c3",  x"6b",  x"c8", -- 14C8
         x"2a",  x"31",  x"01",  x"3e",  x"85",  x"2b",  x"be",  x"20", -- 14D0
         x"fc",  x"c9",  x"cd",  x"82",  x"c8",  x"c0",  x"21",  x"00", -- 14D8
         x"02",  x"36",  x"00",  x"23",  x"36",  x"20",  x"22",  x"33", -- 14E0
         x"01",  x"2a",  x"20",  x"01",  x"22",  x"2f",  x"01",  x"c9", -- 14E8
         x"2a",  x"33",  x"01",  x"c3",  x"50",  x"dd",  x"ed",  x"4b", -- 14F0
         x"39",  x"01",  x"cd",  x"24",  x"d5",  x"2a",  x"20",  x"01", -- 14F8
         x"ed",  x"5b",  x"2f",  x"01",  x"cd",  x"0e",  x"c9",  x"03", -- 1500
         x"2a",  x"31",  x"01",  x"eb",  x"ed",  x"b0",  x"1b",  x"ed", -- 1508
         x"53",  x"33",  x"01",  x"c9",  x"01",  x"28",  x"00",  x"cd", -- 1510
         x"24",  x"d5",  x"3e",  x"0a",  x"cd",  x"40",  x"d8",  x"3e", -- 1518
         x"0b",  x"c3",  x"6b",  x"c8",  x"2a",  x"31",  x"01",  x"11", -- 1520
         x"28",  x"b2",  x"1a",  x"77",  x"23",  x"0b",  x"78",  x"b1", -- 1528
         x"28",  x"0c",  x"1a",  x"b7",  x"13",  x"20",  x"f3",  x"1a", -- 1530
         x"b7",  x"20",  x"f0",  x"2b",  x"18",  x"ed",  x"22",  x"31", -- 1538
         x"01",  x"ed",  x"5b",  x"2f",  x"01",  x"b7",  x"ed",  x"52", -- 1540
         x"d8",  x"ed",  x"53",  x"31",  x"01",  x"cd",  x"c9",  x"c7", -- 1548
         x"21",  x"9c",  x"c1",  x"c3",  x"0b",  x"c8",  x"e5",  x"21", -- 1550
         x"22",  x"01",  x"cb",  x"7e",  x"e1",  x"c9",  x"cd",  x"85", -- 1558
         x"c9",  x"3a",  x"22",  x"01",  x"cb",  x"ff",  x"18",  x"3a", -- 1560
         x"cd",  x"85",  x"c9",  x"cd",  x"e3",  x"d3",  x"ca",  x"1e", -- 1568
         x"d3",  x"2a",  x"27",  x"01",  x"23",  x"3a",  x"22",  x"01", -- 1570
         x"cb",  x"ff",  x"18",  x"2f",  x"cd",  x"c9",  x"c7",  x"21", -- 1578
         x"8f",  x"c2",  x"cd",  x"4a",  x"c9",  x"7c",  x"b7",  x"20", -- 1580
         x"f3",  x"7d",  x"fe",  x"0a",  x"38",  x"ee",  x"32",  x"35", -- 1588
         x"01",  x"cb",  x"3f",  x"cb",  x"3f",  x"cb",  x"3f",  x"06", -- 1590
         x"08",  x"80",  x"32",  x"3b",  x"01",  x"3a",  x"22",  x"01", -- 1598
         x"cb",  x"bf",  x"2a",  x"33",  x"01",  x"22",  x"29",  x"01", -- 15A0
         x"21",  x"01",  x"02",  x"32",  x"22",  x"01",  x"e5",  x"1e", -- 15A8
         x"04",  x"cd",  x"61",  x"d1",  x"e1",  x"3a",  x"35",  x"01", -- 15B0
         x"47",  x"04",  x"e5",  x"7e",  x"b7",  x"28",  x"15",  x"fe", -- 15B8
         x"84",  x"ca",  x"6e",  x"d6",  x"fe",  x"8b",  x"28",  x"31", -- 15C0
         x"fe",  x"89",  x"ca",  x"41",  x"d6",  x"23",  x"10",  x"eb", -- 15C8
         x"2b",  x"c3",  x"a2",  x"d6",  x"cd",  x"56",  x"d5",  x"20", -- 15D0
         x"04",  x"c1",  x"23",  x"18",  x"09",  x"e1",  x"cd",  x"00", -- 15D8
         x"d8",  x"cd",  x"f0",  x"c9",  x"28",  x"0d",  x"e5",  x"ed", -- 15E0
         x"5b",  x"29",  x"01",  x"1b",  x"1b",  x"b7",  x"ed",  x"52", -- 15E8
         x"e1",  x"38",  x"c2",  x"cd",  x"98",  x"c8",  x"c3",  x"5f", -- 15F0
         x"d1",  x"c1",  x"3a",  x"35",  x"01",  x"47",  x"c5",  x"0e", -- 15F8
         x"00",  x"23",  x"e5",  x"7e",  x"23",  x"b7",  x"28",  x"13", -- 1600
         x"0c",  x"10",  x"f8",  x"c1",  x"c1",  x"cd",  x"80",  x"dd", -- 1608
         x"cd",  x"31",  x"c8",  x"c3",  x"b6",  x"d2",  x"2a",  x"25", -- 1610
         x"01",  x"18",  x"f2",  x"cd",  x"56",  x"d5",  x"28",  x"19", -- 1618
         x"e1",  x"f1",  x"91",  x"cb",  x"3f",  x"28",  x"08",  x"47", -- 1620
         x"3e",  x"20",  x"cd",  x"7d",  x"c8",  x"10",  x"fb",  x"7e", -- 1628
         x"23",  x"b7",  x"28",  x"08",  x"cd",  x"7d",  x"c8",  x"18", -- 1630
         x"f6",  x"c1",  x"18",  x"9d",  x"cd",  x"8b",  x"c8",  x"18", -- 1638
         x"a0",  x"e1",  x"3a",  x"35",  x"01",  x"47",  x"0e",  x"01", -- 1640
         x"7e",  x"23",  x"b7",  x"28",  x"ef",  x"fe",  x"89",  x"28", -- 1648
         x"0b",  x"cd",  x"56",  x"d5",  x"c4",  x"7d",  x"c8",  x"0c", -- 1650
         x"10",  x"ee",  x"18",  x"b1",  x"3e",  x"20",  x"cd",  x"56", -- 1658
         x"d5",  x"c4",  x"7d",  x"c8",  x"0c",  x"79",  x"e6",  x"03", -- 1660
         x"28",  x"ee",  x"10",  x"f0",  x"18",  x"9f",  x"3a",  x"35", -- 1668
         x"01",  x"3d",  x"47",  x"e1",  x"7e",  x"23",  x"b7",  x"28", -- 1670
         x"c3",  x"fe",  x"84",  x"28",  x"0a",  x"cd",  x"56",  x"d5", -- 1678
         x"c4",  x"7d",  x"c8",  x"10",  x"ef",  x"18",  x"e5",  x"e5", -- 1680
         x"af",  x"23",  x"be",  x"28",  x"05",  x"10",  x"fa",  x"e1", -- 1688
         x"18",  x"da",  x"cd",  x"56",  x"d5",  x"ca",  x"d9",  x"d5", -- 1690
         x"3e",  x"20",  x"cd",  x"7d",  x"c8",  x"10",  x"fb",  x"e1", -- 1698
         x"18",  x"d2",  x"e5",  x"fe",  x"20",  x"28",  x"43",  x"3a", -- 16A0
         x"3b",  x"01",  x"4f",  x"47",  x"2b",  x"7e",  x"fe",  x"20", -- 16A8
         x"28",  x"38",  x"fe",  x"28",  x"20",  x"03",  x"2b",  x"18", -- 16B0
         x"37",  x"fe",  x"30",  x"38",  x"33",  x"fe",  x"3a",  x"38", -- 16B8
         x"08",  x"fe",  x"40",  x"38",  x"2b",  x"fe",  x"8c",  x"28", -- 16C0
         x"27",  x"10",  x"e1",  x"e1",  x"41",  x"2b",  x"0d",  x"2b", -- 16C8
         x"7e",  x"cb",  x"af",  x"fe",  x"59",  x"28",  x"64",  x"e5", -- 16D0
         x"c5",  x"06",  x"0b",  x"21",  x"35",  x"d8",  x"be",  x"28", -- 16D8
         x"57",  x"23",  x"10",  x"fa",  x"c1",  x"e1",  x"10",  x"e7", -- 16E0
         x"18",  x"50",  x"3e",  x"20",  x"2b",  x"be",  x"28",  x"fa", -- 16E8
         x"c1",  x"d1",  x"cd",  x"dc",  x"d7",  x"cd",  x"56",  x"d5", -- 16F0
         x"ca",  x"c6",  x"d7",  x"21",  x"22",  x"01",  x"cb",  x"6e", -- 16F8
         x"16",  x"19",  x"28",  x"09",  x"cd",  x"f7",  x"d7",  x"cd", -- 1700
         x"00",  x"d8",  x"c3",  x"c6",  x"d7",  x"cd",  x"f7",  x"d7", -- 1708
         x"15",  x"28",  x"f1",  x"7e",  x"fe",  x"20",  x"23",  x"cd", -- 1710
         x"6b",  x"c8",  x"28",  x"f7",  x"7e",  x"b7",  x"28",  x"ed", -- 1718
         x"fe",  x"20",  x"23",  x"cd",  x"6b",  x"c8",  x"20",  x"f4", -- 1720
         x"0d",  x"28",  x"d9",  x"3e",  x"1a",  x"cd",  x"6b",  x"c8", -- 1728
         x"3e",  x"20",  x"cd",  x"6b",  x"c8",  x"23",  x"18",  x"e4", -- 1730
         x"c1",  x"e1",  x"23",  x"d1",  x"cd",  x"dc",  x"d7",  x"e5", -- 1738
         x"ed",  x"5b",  x"a0",  x"b7",  x"3e",  x"8c",  x"cd",  x"6b", -- 1740
         x"c8",  x"0d",  x"28",  x"08",  x"41",  x"7e",  x"cd",  x"6b", -- 1748
         x"c8",  x"23",  x"10",  x"f9",  x"ed",  x"53",  x"a0",  x"b7", -- 1750
         x"e1",  x"cd",  x"31",  x"c8",  x"fe",  x"0d",  x"47",  x"28", -- 1758
         x"34",  x"fe",  x"08",  x"28",  x"0d",  x"fe",  x"09",  x"20", -- 1760
         x"f0",  x"c3",  x"f0",  x"dd",  x"0c",  x"18",  x"ea",  x"23", -- 1768
         x"18",  x"09",  x"3a",  x"3b",  x"01",  x"3d",  x"b9",  x"38", -- 1770
         x"e0",  x"2b",  x"0c",  x"3e",  x"1f",  x"cd",  x"6b",  x"c8", -- 1778
         x"78",  x"cd",  x"6b",  x"c8",  x"3e",  x"1a",  x"cd",  x"6b", -- 1780
         x"c8",  x"3e",  x"8c",  x"cd",  x"6b",  x"c8",  x"3e",  x"08", -- 1788
         x"cd",  x"6b",  x"c8",  x"18",  x"c4",  x"22",  x"25",  x"01", -- 1790
         x"3e",  x"09",  x"cd",  x"6b",  x"c8",  x"41",  x"3e",  x"1f", -- 1798
         x"cd",  x"6b",  x"c8",  x"10",  x"fb",  x"cd",  x"56",  x"d5", -- 17A0
         x"c2",  x"fb",  x"d6",  x"eb",  x"cd",  x"f0",  x"d4",  x"2a", -- 17A8
         x"33",  x"01",  x"e5",  x"03",  x"d1",  x"13",  x"ed",  x"53", -- 17B0
         x"33",  x"01",  x"ed",  x"b8",  x"3e",  x"8c",  x"12",  x"2a", -- 17B8
         x"29",  x"01",  x"23",  x"22",  x"29",  x"01",  x"3a",  x"22", -- 17C0
         x"01",  x"cb",  x"af",  x"fe",  x"52",  x"2a",  x"25",  x"01", -- 17C8
         x"c4",  x"f0",  x"c9",  x"3e",  x"20",  x"23",  x"be",  x"28", -- 17D0
         x"fc",  x"c3",  x"b5",  x"d5",  x"22",  x"25",  x"01",  x"cd", -- 17D8
         x"0e",  x"c9",  x"41",  x"3a",  x"35",  x"01",  x"90",  x"4f", -- 17E0
         x"04",  x"cd",  x"69",  x"c8",  x"eb",  x"c5",  x"7e",  x"cd", -- 17E8
         x"6b",  x"c8",  x"23",  x"10",  x"f9",  x"c1",  x"c9",  x"3e", -- 17F0
         x"10",  x"cd",  x"6b",  x"c8",  x"21",  x"28",  x"b2",  x"c9", -- 17F8
         x"7e",  x"23",  x"b7",  x"ca",  x"8b",  x"c8",  x"fe",  x"8c", -- 1800
         x"20",  x"02",  x"3e",  x"2d",  x"cd",  x"7d",  x"c8",  x"18", -- 1808
         x"ef",  x"4e",  x"cb",  x"d1",  x"54",  x"ce",  x"d1",  x"42", -- 1810
         x"c5",  x"d1",  x"47",  x"a2",  x"d1",  x"4c",  x"a0",  x"d4", -- 1818
         x"57",  x"a5",  x"d4",  x"5a",  x"40",  x"d4",  x"52",  x"7f", -- 1820
         x"d5",  x"46",  x"7e",  x"d1",  x"48",  x"f5",  x"c7",  x"45", -- 1828
         x"5e",  x"d5",  x"03",  x"96",  x"d1",  x"45",  x"41",  x"49", -- 1830
         x"4f",  x"55",  x"80",  x"81",  x"82",  x"86",  x"87",  x"88", -- 1838
         x"cd",  x"4b",  x"d8",  x"21",  x"4f",  x"d8",  x"e5",  x"2a", -- 1840
         x"1e",  x"01",  x"e9",  x"3e",  x"3a",  x"18",  x"02",  x"3e", -- 1848
         x"07",  x"c3",  x"30",  x"dc",  x"c9",  x"a4",  x"e3",  x"88", -- 1850
         x"9e",  x"9b",  x"99",  x"9b",  x"87",  x"99",  x"9c",  x"a5", -- 1858
         x"fb",  x"cb",  x"c0",  x"da",  x"c1",  x"ce",  x"dc",  x"a5", -- 1860
         x"a5",  x"f8",  x"92",  x"f8",  x"c1",  x"cb",  x"c9",  x"a5", -- 1868
         x"ed",  x"92",  x"ed",  x"c4",  x"c1",  x"dc",  x"cd",  x"a5", -- 1870
         x"e3",  x"92",  x"c3",  x"c7",  x"c5",  x"d8",  x"da",  x"c1", -- 1878
         x"c5",  x"c1",  x"cd",  x"da",  x"dc",  x"a5",  x"a5",  x"a8", -- 1880
         x"a5",  x"fb",  x"d8",  x"cd",  x"da",  x"da",  x"db",  x"cb", -- 1888
         x"c0",  x"da",  x"c1",  x"ce",  x"dc",  x"88",  x"98",  x"87", -- 1890
         x"99",  x"a5",  x"a8",  x"a5",  x"f2",  x"cd",  x"c1",  x"c4", -- 1898
         x"cd",  x"c6",  x"c9",  x"ca",  x"db",  x"dc",  x"c9",  x"c6", -- 18A0
         x"cc",  x"88",  x"9a",  x"87",  x"9b",  x"87",  x"9c",  x"a5", -- 18A8
         x"a8",  x"a5",  x"e9",  x"c6",  x"ce",  x"c9",  x"c6",  x"cf", -- 18B0
         x"db",  x"db",  x"d8",  x"c9",  x"cb",  x"cd",  x"a5",  x"a8", -- 18B8
         x"a4",  x"8b",  x"8b",  x"8b",  x"8b",  x"88",  x"e1",  x"e6", -- 18C0
         x"e1",  x"fc",  x"88",  x"8b",  x"8b",  x"8b",  x"8b",  x"a5", -- 18C8
         x"a5",  x"a5",  x"fb",  x"dc",  x"cd",  x"dd",  x"cd",  x"da", -- 18D0
         x"d2",  x"cd",  x"c1",  x"cb",  x"c0",  x"cd",  x"c6",  x"88", -- 18D8
         x"e2",  x"87",  x"e6",  x"a5",  x"a8",  x"a5",  x"88",  x"88", -- 18E0
         x"82",  x"82",  x"88",  x"ec",  x"da",  x"dd",  x"cb",  x"c3", -- 18E8
         x"cd",  x"da",  x"dc",  x"d1",  x"d8",  x"88",  x"82",  x"82", -- 18F0
         x"a5",  x"a5",  x"88",  x"ed",  x"88",  x"92",  x"88",  x"ed", -- 18F8
         x"da",  x"c1",  x"c3",  x"c9",  x"88",  x"fb",  x"88",  x"9e", -- 1900
         x"98",  x"98",  x"9d",  x"a5",  x"88",  x"e3",  x"88",  x"92", -- 1908
         x"88",  x"e3",  x"88",  x"9e",  x"9b",  x"99",  x"9b",  x"87", -- 1910
         x"99",  x"9c",  x"a5",  x"88",  x"e4",  x"88",  x"92",  x"88", -- 1918
         x"e3",  x"88",  x"9e",  x"9b",  x"99",  x"99",  x"87",  x"99", -- 1920
         x"9a",  x"a5",  x"88",  x"e5",  x"88",  x"92",  x"88",  x"e3", -- 1928
         x"88",  x"9e",  x"9b",  x"98",  x"9c",  x"a5",  x"88",  x"fb", -- 1930
         x"88",  x"92",  x"88",  x"fb",  x"88",  x"9e",  x"98",  x"99", -- 1938
         x"98",  x"a5",  x"a5",  x"88",  x"e9",  x"88",  x"92",  x"88", -- 1940
         x"e9",  x"dd",  x"db",  x"cf",  x"c9",  x"ca",  x"cd",  x"88", -- 1948
         x"fe",  x"c1",  x"cc",  x"cd",  x"c7",  x"a5",  x"a5",  x"a8", -- 1950
         x"e1",  x"21",  x"a3",  x"c7",  x"e5",  x"cd",  x"58",  x"c8", -- 1958
         x"21",  x"c0",  x"d8",  x"cd",  x"3d",  x"da",  x"32",  x"19", -- 1960
         x"01",  x"21",  x"e5",  x"d8",  x"cd",  x"0b",  x"c8",  x"11", -- 1968
         x"f1",  x"da",  x"06",  x"06",  x"c3",  x"af",  x"c7",  x"01", -- 1970
         x"0c",  x"02",  x"21",  x"e9",  x"da",  x"ed",  x"b3",  x"01", -- 1978
         x"0a",  x"06",  x"ed",  x"b3",  x"18",  x"11",  x"3a",  x"1c", -- 1980
         x"01",  x"fe",  x"4b",  x"cc",  x"b6",  x"da",  x"cd",  x"98", -- 1988
         x"c8",  x"00",  x"c3",  x"90",  x"dc",  x"00",  x"00",  x"3a", -- 1990
         x"22",  x"01",  x"32",  x"1c",  x"01",  x"c9",  x"c3",  x"c0", -- 1998
         x"dc",  x"cd",  x"7d",  x"c8",  x"c3",  x"07",  x"cc",  x"00", -- 19A0
         x"00",  x"00",  x"00",  x"e1",  x"cd",  x"03",  x"f0",  x"23", -- 19A8
         x"08",  x"4d",  x"6f",  x"64",  x"75",  x"6c",  x"2d",  x"45", -- 19B0
         x"72",  x"72",  x"6f",  x"72",  x"00",  x"cd",  x"03",  x"f0", -- 19B8
         x"0e",  x"c9",  x"cd",  x"9e",  x"d9",  x"21",  x"62",  x"da", -- 19C0
         x"22",  x"be",  x"b7",  x"21",  x"55",  x"d8",  x"cd",  x"3d", -- 19C8
         x"da",  x"f5",  x"21",  x"88",  x"d8",  x"cd",  x"3d",  x"da", -- 19D0
         x"d6",  x"10",  x"f5",  x"21",  x"9b",  x"d8",  x"cd",  x"3d", -- 19D8
         x"da",  x"f5",  x"21",  x"b1",  x"d8",  x"cd",  x"43",  x"da", -- 19E0
         x"22",  x"1a",  x"01",  x"cd",  x"b6",  x"da",  x"cd",  x"c0", -- 19E8
         x"da",  x"3e",  x"41",  x"cd",  x"c2",  x"da",  x"f1",  x"d6", -- 19F0
         x"10",  x"87",  x"87",  x"3c",  x"cd",  x"bd",  x"da",  x"3e", -- 19F8
         x"57",  x"cd",  x"c2",  x"da",  x"f1",  x"fe",  x"01",  x"28", -- 1A00
         x"01",  x"af",  x"cd",  x"bd",  x"da",  x"f1",  x"fe",  x"50", -- 1A08
         x"28",  x"0a",  x"fe",  x"4b",  x"20",  x"04",  x"3e",  x"0f", -- 1A10
         x"18",  x"02",  x"3e",  x"4d",  x"cd",  x"bd",  x"da",  x"3e", -- 1A18
         x"52",  x"cd",  x"c2",  x"da",  x"3e",  x"02",  x"cd",  x"c2", -- 1A20
         x"da",  x"3e",  x"0d",  x"18",  x"50",  x"3e",  x"01",  x"32", -- 1A28
         x"1a",  x"01",  x"cd",  x"9e",  x"d9",  x"21",  x"54",  x"da", -- 1A30
         x"22",  x"be",  x"b7",  x"18",  x"ec",  x"cd",  x"29",  x"c8", -- 1A38
         x"cb",  x"af",  x"c9",  x"cd",  x"0b",  x"c8",  x"cd",  x"03", -- 1A40
         x"f0",  x"17",  x"cd",  x"03",  x"f0",  x"22",  x"2a",  x"82", -- 1A48
         x"b7",  x"c3",  x"e4",  x"c8",  x"c3",  x"5d",  x"db",  x"cb", -- 1A50
         x"7f",  x"28",  x"22",  x"e5",  x"c5",  x"21",  x"e0",  x"da", -- 1A58
         x"18",  x"0c",  x"c3",  x"84",  x"db",  x"cb",  x"7f",  x"28", -- 1A60
         x"14",  x"e5",  x"c5",  x"21",  x"d7",  x"da",  x"d6",  x"80", -- 1A68
         x"fe",  x"09",  x"38",  x"02",  x"3e",  x"04",  x"4f",  x"06", -- 1A70
         x"00",  x"09",  x"7e",  x"c1",  x"e1",  x"c3",  x"08",  x"de", -- 1A78
         x"00",  x"32",  x"1d",  x"01",  x"c9",  x"c3",  x"00",  x"df", -- 1A80
         x"00",  x"b7",  x"28",  x"17",  x"f1",  x"fe",  x"0d",  x"c8", -- 1A88
         x"fe",  x"0a",  x"20",  x"03",  x"af",  x"18",  x"ea",  x"c3", -- 1A90
         x"18",  x"de",  x"3a",  x"19",  x"01",  x"fe",  x"4a",  x"28", -- 1A98
         x"02",  x"f1",  x"c9",  x"f1",  x"cd",  x"c2",  x"da",  x"fe", -- 1AA0
         x"0d",  x"c0",  x"3a",  x"1a",  x"01",  x"c3",  x"10",  x"dc", -- 1AA8
         x"cd",  x"c2",  x"da",  x"10",  x"fb",  x"c9",  x"cd",  x"c0", -- 1AB0
         x"da",  x"3e",  x"40",  x"18",  x"05",  x"cd",  x"c2",  x"da", -- 1AB8
         x"3e",  x"1b",  x"c5",  x"f5",  x"db",  x"0a",  x"cb",  x"57", -- 1AC0
         x"20",  x"08",  x"3e",  x"01",  x"cd",  x"03",  x"f0",  x"14", -- 1AC8
         x"18",  x"f2",  x"f1",  x"d3",  x"08",  x"c1",  x"c9",  x"7b", -- 1AD0
         x"7c",  x"7d",  x"7e",  x"20",  x"20",  x"5b",  x"5c",  x"5d", -- 1AD8
         x"7b",  x"7c",  x"7d",  x"83",  x"20",  x"20",  x"5b",  x"5c", -- 1AE0
         x"5d",  x"47",  x"5b",  x"04",  x"04",  x"03",  x"20",  x"05", -- 1AE8
         x"6a",  x"45",  x"2d",  x"da",  x"4b",  x"c2",  x"d9",  x"41", -- 1AF0
         x"86",  x"d9",  x"4c",  x"48",  x"db",  x"4d",  x"40",  x"dc", -- 1AF8
         x"53",  x"03",  x"db",  x"3e",  x"01",  x"32",  x"1a",  x"01", -- 1B00
         x"cd",  x"9e",  x"d9",  x"21",  x"11",  x"db",  x"c3",  x"38", -- 1B08
         x"da",  x"cd",  x"6b",  x"c8",  x"cb",  x"7f",  x"ca",  x"7d", -- 1B10
         x"da",  x"e5",  x"c5",  x"21",  x"21",  x"db",  x"c3",  x"6e", -- 1B18
         x"da",  x"84",  x"94",  x"81",  x"e1",  x"20",  x"20",  x"8e", -- 1B20
         x"99",  x"9a",  x"07",  x"59",  x"04",  x"04",  x"03",  x"20", -- 1B28
         x"05",  x"6a",  x"1b",  x"5b",  x"31",  x"34",  x"34",  x"7d", -- 1B30
         x"1b",  x"5b",  x"31",  x"32",  x"30",  x"7a",  x"1b",  x"52", -- 1B38
         x"02",  x"00",  x"1b",  x"5b",  x"30",  x"20",  x"4b",  x"0a", -- 1B40
         x"c3",  x"80",  x"dc",  x"01",  x"0c",  x"02",  x"21",  x"2a", -- 1B48
         x"db",  x"cd",  x"7d",  x"d9",  x"21",  x"ea",  x"db",  x"cd", -- 1B50
         x"3d",  x"da",  x"f5",  x"18",  x"10",  x"cd",  x"6b",  x"c8", -- 1B58
         x"fe",  x"87",  x"c2",  x"57",  x"da",  x"3e",  x"5c",  x"c3", -- 1B60
         x"a4",  x"da",  x"ff",  x"ff",  x"ff",  x"21",  x"b1",  x"d8", -- 1B68
         x"cd",  x"43",  x"da",  x"22",  x"1a",  x"01",  x"06",  x"16", -- 1B70
         x"21",  x"32",  x"db",  x"7e",  x"cd",  x"c2",  x"da",  x"23", -- 1B78
         x"10",  x"f9",  x"18",  x"1e",  x"cd",  x"6b",  x"c8",  x"fe", -- 1B80
         x"87",  x"c2",  x"65",  x"da",  x"c3",  x"65",  x"db",  x"cd", -- 1B88
         x"6b",  x"c8",  x"fe",  x"87",  x"c2",  x"51",  x"dc",  x"c3", -- 1B90
         x"65",  x"db",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1B98
         x"ff",  x"ff",  x"f1",  x"fe",  x"12",  x"20",  x"08",  x"cd", -- 1BA0
         x"be",  x"db",  x"3e",  x"32",  x"cd",  x"c8",  x"db",  x"fe", -- 1BA8
         x"15",  x"20",  x"08",  x"cd",  x"be",  x"db",  x"3e",  x"33", -- 1BB0
         x"cd",  x"c8",  x"db",  x"c3",  x"29",  x"da",  x"3e",  x"1b", -- 1BB8
         x"cd",  x"c2",  x"da",  x"3e",  x"5b",  x"c3",  x"c2",  x"da", -- 1BC0
         x"cd",  x"c2",  x"da",  x"3e",  x"20",  x"cd",  x"c2",  x"da", -- 1BC8
         x"3e",  x"4b",  x"c3",  x"c2",  x"da",  x"a5",  x"fb",  x"cb", -- 1BD0
         x"c0",  x"da",  x"c9",  x"cd",  x"cf",  x"db",  x"cb",  x"c0", -- 1BD8
         x"da",  x"c1",  x"ce",  x"dc",  x"88",  x"98",  x"87",  x"99", -- 1BE0
         x"a5",  x"a8",  x"a4",  x"e3",  x"88",  x"9e",  x"9b",  x"99", -- 1BE8
         x"99",  x"87",  x"99",  x"9a",  x"a5",  x"a5",  x"fb",  x"cb", -- 1BF0
         x"c0",  x"da",  x"c1",  x"ce",  x"dc",  x"ca",  x"da",  x"cd", -- 1BF8
         x"c1",  x"dc",  x"cd",  x"88",  x"98",  x"84",  x"9a",  x"84", -- 1C00
         x"9d",  x"a5",  x"a8",  x"c9",  x"f1",  x"c3",  x"98",  x"da", -- 1C08
         x"c5",  x"47",  x"3e",  x"20",  x"cd",  x"c2",  x"da",  x"10", -- 1C10
         x"fb",  x"c1",  x"c9",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C18
         x"cd",  x"58",  x"c8",  x"21",  x"c0",  x"d8",  x"cd",  x"35", -- 1C20
         x"da",  x"32",  x"18",  x"01",  x"c9",  x"00",  x"00",  x"00", -- 1C28
         x"32",  x"a3",  x"b7",  x"2a",  x"1e",  x"01",  x"22",  x"a4", -- 1C30
         x"b7",  x"c9",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C38
         x"3e",  x"01",  x"32",  x"1a",  x"01",  x"cd",  x"9e",  x"d9", -- 1C40
         x"21",  x"4e",  x"dc",  x"c3",  x"38",  x"da",  x"c3",  x"8f", -- 1C48
         x"db",  x"cb",  x"7f",  x"ca",  x"7d",  x"da",  x"e5",  x"c5", -- 1C50
         x"21",  x"5e",  x"dc",  x"c3",  x"6e",  x"da",  x"7b",  x"7c", -- 1C58
         x"7d",  x"7e",  x"20",  x"20",  x"5b",  x"5c",  x"5d",  x"00", -- 1C60
         x"ff",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1C68
         x"3a",  x"22",  x"01",  x"cb",  x"af",  x"fe",  x"4c",  x"c2", -- 1C70
         x"77",  x"d9",  x"c9",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C78
         x"cd",  x"9e",  x"d9",  x"21",  x"62",  x"da",  x"22",  x"be", -- 1C80
         x"b7",  x"c3",  x"4b",  x"db",  x"ff",  x"ff",  x"ff",  x"ff", -- 1C88
         x"e5",  x"d5",  x"16",  x"3e",  x"3e",  x"01",  x"2e",  x"08", -- 1C90
         x"d5",  x"f5",  x"cd",  x"03",  x"f0",  x"26",  x"7c",  x"fe", -- 1C98
         x"ee",  x"28",  x"0e",  x"7d",  x"c6",  x"04",  x"6f",  x"f1", -- 1CA0
         x"d1",  x"15",  x"20",  x"ec",  x"d1",  x"e1",  x"c3",  x"97", -- 1CA8
         x"d9",  x"f1",  x"d1",  x"3c",  x"16",  x"00",  x"5a",  x"cd", -- 1CB0
         x"03",  x"f0",  x"26",  x"18",  x"ef",  x"00",  x"00",  x"00", -- 1CB8
         x"e5",  x"d5",  x"16",  x"3e",  x"3e",  x"01",  x"2e",  x"08", -- 1CC0
         x"d5",  x"f5",  x"cd",  x"03",  x"f0",  x"26",  x"7c",  x"fe", -- 1CC8
         x"ee",  x"28",  x"0e",  x"7d",  x"c6",  x"04",  x"6f",  x"f1", -- 1CD0
         x"d1",  x"15",  x"20",  x"ec",  x"d1",  x"e1",  x"c3",  x"ab", -- 1CD8
         x"d9",  x"f1",  x"d1",  x"3c",  x"16",  x"01",  x"5a",  x"cd", -- 1CE0
         x"03",  x"f0",  x"26",  x"d1",  x"e1",  x"c3",  x"70",  x"dc", -- 1CE8
         x"cd",  x"0b",  x"c8",  x"21",  x"4b",  x"45",  x"22",  x"00", -- 1CF0
         x"b7",  x"21",  x"59",  x"01",  x"22",  x"02",  x"b7",  x"af", -- 1CF8
         x"3e",  x"7f",  x"01",  x"00",  x"20",  x"11",  x"00",  x"b7", -- 1D00
         x"21",  x"00",  x"e0",  x"cd",  x"03",  x"f0",  x"1d",  x"26", -- 1D08
         x"e6",  x"38",  x"15",  x"2e",  x"00",  x"22",  x"a8",  x"b7", -- 1D10
         x"22",  x"ac",  x"b7",  x"06",  x"04",  x"21",  x"00",  x"b7", -- 1D18
         x"36",  x"00",  x"23",  x"10",  x"fb",  x"c3",  x"dd",  x"c7", -- 1D20
         x"26",  x"fe",  x"18",  x"e7",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D28
         x"cd",  x"5a",  x"d1",  x"cd",  x"69",  x"c8",  x"c3",  x"4e", -- 1D30
         x"d1",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D38
         x"e1",  x"c3",  x"a3",  x"c7",  x"ff",  x"cd",  x"03",  x"f0", -- 1D40
         x"23",  x"0b",  x"00",  x"c9",  x"ff",  x"ff",  x"ff",  x"ff", -- 1D48
         x"b7",  x"ed",  x"52",  x"44",  x"4d",  x"f5",  x"78",  x"b1", -- 1D50
         x"20",  x"01",  x"03",  x"f1",  x"c9",  x"ff",  x"ff",  x"ff", -- 1D58
         x"1e",  x"05",  x"2e",  x"07",  x"cd",  x"4e",  x"c8",  x"11", -- 1D60
         x"da",  x"ca",  x"c3",  x"a0",  x"ca",  x"ff",  x"ff",  x"ff", -- 1D68
         x"e1",  x"eb",  x"ed",  x"b0",  x"eb",  x"22",  x"33",  x"01", -- 1D70
         x"2b",  x"2b",  x"c3",  x"d8",  x"dd",  x"ff",  x"ff",  x"ff", -- 1D78
         x"cd",  x"03",  x"f0",  x"23",  x"0a",  x"0d",  x"00",  x"cd", -- 1D80
         x"03",  x"f0",  x"19",  x"cd",  x"03",  x"f0",  x"23",  x"0a", -- 1D88
         x"00",  x"00",  x"c3",  x"c9",  x"c7",  x"ff",  x"ff",  x"ff", -- 1D90
         x"cd",  x"03",  x"f0",  x"23",  x"08",  x"00",  x"21",  x"5c", -- 1D98
         x"c1",  x"c3",  x"29",  x"cb",  x"ff",  x"ff",  x"ff",  x"ff", -- 1DA0
         x"1e",  x"06",  x"2e",  x"00",  x"cd",  x"4e",  x"c8",  x"11", -- 1DA8
         x"a0",  x"c8",  x"c3",  x"ad",  x"c7",  x"ff",  x"ff",  x"ff", -- 1DB0
         x"1e",  x"04",  x"2e",  x"07",  x"cd",  x"4e",  x"c8",  x"11", -- 1DB8
         x"56",  x"cf",  x"c3",  x"53",  x"cf",  x"ff",  x"ff",  x"ff", -- 1DC0
         x"1e",  x"07",  x"2e",  x"00",  x"cd",  x"4e",  x"c8",  x"21", -- 1DC8
         x"4b",  x"c1",  x"c3",  x"17",  x"d1",  x"ff",  x"ff",  x"ff", -- 1DD0
         x"23",  x"cd",  x"0b",  x"c9",  x"eb",  x"af",  x"57",  x"5f", -- 1DD8
         x"ed",  x"b1",  x"20",  x"03",  x"13",  x"18",  x"f9",  x"13", -- 1DE0
         x"ed",  x"53",  x"37",  x"01",  x"c9",  x"ff",  x"ff",  x"ff", -- 1DE8
         x"fe",  x"09",  x"c2",  x"59",  x"d7",  x"79",  x"fe",  x"00", -- 1DF0
         x"ca",  x"59",  x"d7",  x"0d",  x"c2",  x"6f",  x"d7",  x"c3", -- 1DF8
         x"6c",  x"d7",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1E00
         x"fe",  x"5e",  x"ca",  x"81",  x"da",  x"fe",  x"5f",  x"c2", -- 1E08
         x"85",  x"da",  x"c3",  x"81",  x"da",  x"ff",  x"ff",  x"ff", -- 1E10
         x"f5",  x"3a",  x"1d",  x"01",  x"fe",  x"5e",  x"20",  x"07", -- 1E18
         x"f1",  x"d6",  x"20",  x"f5",  x"c3",  x"9a",  x"da",  x"f1", -- 1E20
         x"18",  x"f9",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1E28
         x"cd",  x"03",  x"f0",  x"23",  x"0a",  x"0d",  x"61",  x"6c", -- 1E30
         x"74",  x"65",  x"72",  x"20",  x"54",  x"61",  x"62",  x"75", -- 1E38
         x"6c",  x"61",  x"74",  x"6f",  x"72",  x"3a",  x"0a",  x"0d", -- 1E40
         x"00",  x"3a",  x"00",  x"01",  x"cd",  x"03",  x"f0",  x"1c", -- 1E48
         x"cd",  x"03",  x"f0",  x"2c",  x"cd",  x"03",  x"f0",  x"23", -- 1E50
         x"6e",  x"65",  x"75",  x"65",  x"72",  x"20",  x"54",  x"61", -- 1E58
         x"62",  x"75",  x"6c",  x"61",  x"74",  x"6f",  x"72",  x"3a", -- 1E60
         x"0a",  x"0d",  x"00",  x"cd",  x"03",  x"f0",  x"17",  x"cd", -- 1E68
         x"03",  x"f0",  x"18",  x"30",  x"09",  x"cd",  x"03",  x"f0", -- 1E70
         x"23",  x"0b",  x"0b",  x"00",  x"18",  x"d6",  x"3a",  x"97", -- 1E78
         x"b7",  x"b7",  x"28",  x"09",  x"fe",  x"0a",  x"30",  x"ed", -- 1E80
         x"00",  x"00",  x"32",  x"00",  x"01",  x"c9",  x"ff",  x"ff", -- 1E88
         x"cd",  x"31",  x"c8",  x"fe",  x"18",  x"28",  x"03",  x"c3", -- 1E90
         x"33",  x"d2",  x"2a",  x"a0",  x"b7",  x"e5",  x"3a",  x"00", -- 1E98
         x"01",  x"47",  x"af",  x"80",  x"bd",  x"38",  x"fc",  x"20", -- 1EA0
         x"01",  x"80",  x"fe",  x"28",  x"30",  x"0e",  x"f5",  x"47", -- 1EA8
         x"cd",  x"d8",  x"de",  x"f1",  x"e1",  x"6f",  x"22",  x"a0", -- 1EB0
         x"b7",  x"c3",  x"30",  x"d2",  x"06",  x"28",  x"cd",  x"d8", -- 1EB8
         x"de",  x"e1",  x"2e",  x"00",  x"3a",  x"a1",  x"b7",  x"3c", -- 1EC0
         x"47",  x"3a",  x"9f",  x"b7",  x"90",  x"28",  x"06",  x"24", -- 1EC8
         x"22",  x"a0",  x"b7",  x"18",  x"e4",  x"c3",  x"d8",  x"d2", -- 1ED0
         x"d5",  x"2a",  x"a0",  x"b7",  x"2e",  x"00",  x"22",  x"a0", -- 1ED8
         x"b7",  x"2a",  x"a0",  x"b7",  x"e5",  x"d1",  x"c5",  x"cd", -- 1EE0
         x"03",  x"f0",  x"32",  x"c1",  x"7e",  x"fe",  x"00",  x"20", -- 1EE8
         x"02",  x"3e",  x"20",  x"cd",  x"03",  x"f0",  x"24",  x"10", -- 1EF0
         x"e8",  x"d1",  x"c9",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1EF8
         x"f5",  x"fe",  x"5c",  x"20",  x"06",  x"32",  x"01",  x"01", -- 1F00
         x"c3",  x"a1",  x"da",  x"fe",  x"0a",  x"20",  x"17",  x"3a", -- 1F08
         x"01",  x"01",  x"fe",  x"5c",  x"20",  x"06",  x"af",  x"32", -- 1F10
         x"01",  x"01",  x"f1",  x"c9",  x"3a",  x"1d",  x"01",  x"b7", -- 1F18
         x"ca",  x"a3",  x"da",  x"c3",  x"8c",  x"da",  x"3a",  x"01", -- 1F20
         x"01",  x"fe",  x"5c",  x"20",  x"ef",  x"18",  x"eb",  x"cd", -- 1F28
         x"0b",  x"c8",  x"21",  x"02",  x"01",  x"36",  x"00",  x"23", -- 1F30
         x"36",  x"00",  x"2a",  x"33",  x"01",  x"e5",  x"11",  x"01", -- 1F38
         x"02",  x"af",  x"ed",  x"52",  x"20",  x"19",  x"e5",  x"21", -- 1F40
         x"1a",  x"01",  x"22",  x"a0",  x"b7",  x"e1",  x"cd",  x"14", -- 1F48
         x"c9",  x"e1",  x"21",  x"b6",  x"c2",  x"cd",  x"0b",  x"c8", -- 1F50
         x"21",  x"00",  x"05",  x"22",  x"a0",  x"b7",  x"c9",  x"e1", -- 1F58
         x"2b",  x"e5",  x"af",  x"ed",  x"52",  x"28",  x"df",  x"44", -- 1F60
         x"4d",  x"e1",  x"eb",  x"57",  x"5f",  x"7e",  x"fe",  x"5c", -- 1F68
         x"28",  x"0f",  x"fe",  x"5e",  x"28",  x"14",  x"b7",  x"28", -- 1F70
         x"22",  x"23",  x"0b",  x"78",  x"b1",  x"20",  x"ee",  x"18", -- 1F78
         x"1d",  x"3a",  x"02",  x"01",  x"3c",  x"32",  x"02",  x"01", -- 1F80
         x"18",  x"07",  x"3a",  x"03",  x"01",  x"3c",  x"32",  x"03", -- 1F88
         x"01",  x"23",  x"0b",  x"78",  x"b1",  x"28",  x"07",  x"7e", -- 1F90
         x"b7",  x"20",  x"f6",  x"13",  x"18",  x"db",  x"21",  x"1a", -- 1F98
         x"01",  x"22",  x"a0",  x"b7",  x"e5",  x"eb",  x"cd",  x"14", -- 1FA0
         x"c9",  x"21",  x"b6",  x"c2",  x"cd",  x"0b",  x"c8",  x"e1", -- 1FA8
         x"24",  x"22",  x"a0",  x"b7",  x"cd",  x"03",  x"f0",  x"23", -- 1FB0
         x"64",  x"61",  x"76",  x"6f",  x"6e",  x"3a",  x"00",  x"24", -- 1FB8
         x"22",  x"a0",  x"b7",  x"e5",  x"3a",  x"02",  x"01",  x"26", -- 1FC0
         x"00",  x"6f",  x"cd",  x"14",  x"c9",  x"cd",  x"03",  x"f0", -- 1FC8
         x"23",  x"52",  x"2d",  x"5a",  x"65",  x"69",  x"6c",  x"65", -- 1FD0
         x"6e",  x"00",  x"e1",  x"24",  x"22",  x"a0",  x"b7",  x"3a", -- 1FD8
         x"03",  x"01",  x"26",  x"00",  x"6f",  x"cd",  x"14",  x"c9", -- 1FE0
         x"cd",  x"03",  x"f0",  x"23",  x"53",  x"2d",  x"5a",  x"65", -- 1FE8
         x"69",  x"6c",  x"65",  x"6e",  x"00",  x"c3",  x"58",  x"df", -- 1FF0
         x"79",  x"f8",  x"6a",  x"31",  x"50",  x"9d",  x"e3",  x"75"  -- 1FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
