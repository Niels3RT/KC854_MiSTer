library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity caos_c is
    generic(
        ADDR_WIDTH   : integer := 12
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end caos_c;

architecture rtl of caos_c is
    type rom4096x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom4096x8 := (
         x"d5",  x"2e",  x"08",  x"e5",  x"3e",  x"01",  x"cd",  x"04", -- 0000
         x"e4",  x"7c",  x"3c",  x"28",  x"0f",  x"7d",  x"cd",  x"59", -- 0008
         x"f3",  x"7c",  x"cd",  x"59",  x"f3",  x"7a",  x"cd",  x"76", -- 0010
         x"f3",  x"cd",  x"6b",  x"f3",  x"e1",  x"7d",  x"c6",  x"04", -- 0018
         x"6f",  x"30",  x"e0",  x"cd",  x"6b",  x"f3",  x"d1",  x"c9", -- 0020
         x"d5",  x"cd",  x"ee",  x"f1",  x"43",  x"41",  x"4f",  x"53", -- 0028
         x"00",  x"3e",  x"45",  x"cd",  x"29",  x"e3",  x"db",  x"88", -- 0030
         x"0f",  x"38",  x"05",  x"cd",  x"ec",  x"c0",  x"18",  x"03", -- 0038
         x"cd",  x"e2",  x"c0",  x"cd",  x"ee",  x"f1",  x"52",  x"4f", -- 0040
         x"4d",  x"43",  x"20",  x"00",  x"dd",  x"7e",  x"04",  x"cb", -- 0048
         x"3f",  x"cb",  x"3f",  x"cb",  x"3f",  x"cb",  x"3f",  x"cb", -- 0050
         x"3f",  x"2f",  x"e6",  x"33",  x"cd",  x"29",  x"e3",  x"db", -- 0058
         x"88",  x"5f",  x"07",  x"38",  x"05",  x"cd",  x"ec",  x"c0", -- 0060
         x"18",  x"03",  x"cd",  x"e2",  x"c0",  x"cd",  x"da",  x"c0", -- 0068
         x"3e",  x"30",  x"cd",  x"29",  x"e3",  x"cb",  x"4b",  x"20", -- 0070
         x"05",  x"cd",  x"ec",  x"c0",  x"18",  x"03",  x"cd",  x"e2", -- 0078
         x"c0",  x"cd",  x"da",  x"c0",  x"3e",  x"34",  x"cd",  x"29", -- 0080
         x"e3",  x"dd",  x"cb",  x"04",  x"46",  x"20",  x"05",  x"cd", -- 0088
         x"ec",  x"c0",  x"18",  x"03",  x"cd",  x"e2",  x"c0",  x"cd", -- 0090
         x"da",  x"c0",  x"cd",  x"ee",  x"f1",  x"38",  x"20",  x"00", -- 0098
         x"dd",  x"7e",  x"01",  x"cb",  x"3f",  x"cb",  x"3f",  x"cb", -- 00A0
         x"3f",  x"cb",  x"3f",  x"c6",  x"2e",  x"cd",  x"29",  x"e3", -- 00A8
         x"db",  x"89",  x"cb",  x"6f",  x"20",  x"05",  x"cd",  x"ec", -- 00B0
         x"c0",  x"18",  x"03",  x"cd",  x"e2",  x"c0",  x"dd",  x"7e", -- 00B8
         x"01",  x"5f",  x"cd",  x"ee",  x"f1",  x"42",  x"49",  x"4c", -- 00C0
         x"44",  x"20",  x"00",  x"cb",  x"53",  x"3e",  x"30",  x"28", -- 00C8
         x"01",  x"3c",  x"cd",  x"29",  x"e3",  x"cd",  x"6b",  x"f3", -- 00D0
         x"d1",  x"c9",  x"cd",  x"ee",  x"f1",  x"52",  x"41",  x"4d", -- 00D8
         x"00",  x"c9",  x"cd",  x"ee",  x"f1",  x"20",  x"4f",  x"4e", -- 00E0
         x"0d",  x"0a",  x"00",  x"c9",  x"cd",  x"ee",  x"f1",  x"20", -- 00E8
         x"4f",  x"46",  x"46",  x"0d",  x"0a",  x"00",  x"c9",  x"21", -- 00F0
         x"00",  x"b9",  x"01",  x"f0",  x"0c",  x"0c",  x"79",  x"cd", -- 00F8
         x"eb",  x"f1",  x"20",  x"3a",  x"00",  x"cd",  x"cf",  x"f6", -- 0100
         x"cd",  x"6b",  x"f3",  x"10",  x"f0",  x"c9",  x"af",  x"3e", -- 0108
         x"ff",  x"5f",  x"57",  x"3c",  x"13",  x"13",  x"ed",  x"52", -- 0110
         x"f2",  x"13",  x"c1",  x"c9",  x"06",  x"00",  x"1e",  x"09", -- 0118
         x"7a",  x"1f",  x"1d",  x"c8",  x"57",  x"78",  x"30",  x"01", -- 0120
         x"81",  x"1f",  x"47",  x"18",  x"f3",  x"f5",  x"fe",  x"0a", -- 0128
         x"30",  x"2e",  x"7a",  x"a7",  x"28",  x"2a",  x"84",  x"38", -- 0130
         x"27",  x"fe",  x"21",  x"30",  x"23",  x"7b",  x"a7",  x"28", -- 0138
         x"1f",  x"85",  x"38",  x"1c",  x"fe",  x"29",  x"30",  x"18", -- 0140
         x"f1",  x"d5",  x"e5",  x"cd",  x"bb",  x"f6",  x"e1",  x"d1", -- 0148
         x"22",  x"9c",  x"b7",  x"ed",  x"53",  x"9e",  x"b7",  x"ed", -- 0150
         x"43",  x"a0",  x"b7",  x"32",  x"9b",  x"b7",  x"a7",  x"c9", -- 0158
         x"f1",  x"37",  x"c9",  x"3e",  x"1f",  x"a5",  x"17",  x"17", -- 0160
         x"17",  x"6f",  x"3a",  x"81",  x"b7",  x"fe",  x"02",  x"7b", -- 0168
         x"30",  x"03",  x"3a",  x"a3",  x"b7",  x"e6",  x"07",  x"b5", -- 0170
         x"32",  x"a3",  x"b7",  x"c9",  x"2a",  x"84",  x"b7",  x"ed", -- 0178
         x"5b",  x"88",  x"b7",  x"d9",  x"2a",  x"82",  x"b7",  x"ed", -- 0180
         x"5b",  x"86",  x"b7",  x"af",  x"ed",  x"52",  x"30",  x"07", -- 0188
         x"19",  x"eb",  x"d9",  x"eb",  x"d9",  x"18",  x"f4",  x"d9", -- 0190
         x"d5",  x"ed",  x"52",  x"30",  x"06",  x"19",  x"eb",  x"f6", -- 0198
         x"01",  x"18",  x"f6",  x"e5",  x"d9",  x"c1",  x"e5",  x"ed", -- 01A0
         x"42",  x"e1",  x"c5",  x"30",  x"03",  x"e3",  x"f6",  x"02", -- 01A8
         x"e5",  x"44",  x"4d",  x"d9",  x"c1",  x"d1",  x"60",  x"69", -- 01B0
         x"cb",  x"3c",  x"cb",  x"1d",  x"d9",  x"e1",  x"eb",  x"cd", -- 01B8
         x"e8",  x"f7",  x"d9",  x"a7",  x"ed",  x"52",  x"30",  x"01", -- 01C0
         x"09",  x"d9",  x"cb",  x"4f",  x"20",  x"04",  x"23",  x"30", -- 01C8
         x"0b",  x"a7",  x"cb",  x"47",  x"13",  x"28",  x"02",  x"1b", -- 01D0
         x"1b",  x"30",  x"01",  x"23",  x"08",  x"78",  x"b1",  x"c8", -- 01D8
         x"0b",  x"08",  x"18",  x"db",  x"e5",  x"d5",  x"c5",  x"2a", -- 01E0
         x"d3",  x"b7",  x"7d",  x"e6",  x"07",  x"cb",  x"3c",  x"cb", -- 01E8
         x"1d",  x"cb",  x"3c",  x"cb",  x"1d",  x"cb",  x"3c",  x"cb", -- 01F0
         x"1d",  x"c6",  x"f8",  x"4f",  x"06",  x"fd",  x"3a",  x"d5", -- 01F8
         x"b7",  x"2f",  x"67",  x"0a",  x"cd",  x"4e",  x"e0",  x"38", -- 0200
         x"16",  x"47",  x"4e",  x"2f",  x"a1",  x"77",  x"dd",  x"7e", -- 0208
         x"01",  x"5f",  x"ee",  x"02",  x"f3",  x"d3",  x"84",  x"56", -- 0210
         x"7b",  x"d3",  x"84",  x"fb",  x"78",  x"a1",  x"7a",  x"c1", -- 0218
         x"d1",  x"e1",  x"c9",  x"cd",  x"54",  x"f3",  x"e5",  x"41", -- 0220
         x"cd",  x"4a",  x"f6",  x"23",  x"cd",  x"59",  x"f3",  x"10", -- 0228
         x"f7",  x"e1",  x"41",  x"3e",  x"09",  x"cd",  x"1d",  x"f2", -- 0230
         x"cd",  x"4a",  x"f6",  x"23",  x"cd",  x"2a",  x"f6",  x"10", -- 0238
         x"f7",  x"c9",  x"fe",  x"03",  x"30",  x"08",  x"0e",  x"08", -- 0240
         x"fe",  x"02",  x"30",  x"02",  x"1e",  x"04",  x"d5",  x"cd", -- 0248
         x"23",  x"c2",  x"cd",  x"6b",  x"f3",  x"cd",  x"de",  x"e3", -- 0250
         x"38",  x"06",  x"1d",  x"20",  x"f2",  x"cd",  x"17",  x"f2", -- 0258
         x"d1",  x"fe",  x"03",  x"c8",  x"fe",  x"13",  x"20",  x"e6", -- 0260
         x"18",  x"02",  x"0e",  x"01",  x"cd",  x"23",  x"c2",  x"3e", -- 0268
         x"05",  x"32",  x"a0",  x"b7",  x"cd",  x"34",  x"f3",  x"e5", -- 0270
         x"cd",  x"92",  x"f3",  x"7e",  x"e1",  x"38",  x"51",  x"a7", -- 0278
         x"28",  x"ea",  x"2a",  x"97",  x"b7",  x"e5",  x"cd",  x"92", -- 0280
         x"f3",  x"7e",  x"a7",  x"23",  x"7e",  x"e1",  x"28",  x"04", -- 0288
         x"cd",  x"62",  x"f6",  x"23",  x"1a",  x"fe",  x"2e",  x"c8", -- 0290
         x"fe",  x"2c",  x"20",  x"05",  x"13",  x"1a",  x"13",  x"18", -- 0298
         x"ef",  x"fe",  x"3a",  x"20",  x"03",  x"2b",  x"18",  x"c4", -- 02A0
         x"fe",  x"2f",  x"20",  x"0b",  x"13",  x"cd",  x"92",  x"f3", -- 02A8
         x"38",  x"1e",  x"2a",  x"97",  x"b7",  x"18",  x"b5",  x"fe", -- 02B0
         x"27",  x"20",  x"0e",  x"13",  x"1a",  x"13",  x"a7",  x"28", -- 02B8
         x"ab",  x"fe",  x"27",  x"28",  x"cf",  x"77",  x"23",  x"18", -- 02C0
         x"f3",  x"a7",  x"28",  x"a0",  x"fe",  x"20",  x"28",  x"b5", -- 02C8
         x"cd",  x"61",  x"f3",  x"18",  x"97",  x"21",  x"81",  x"b7", -- 02D0
         x"7e",  x"fe",  x"03",  x"30",  x"24",  x"06",  x"08",  x"cd", -- 02D8
         x"b1",  x"c3",  x"38",  x"56",  x"21",  x"e2",  x"f9",  x"22", -- 02E0
         x"99",  x"b7",  x"11",  x"06",  x"fa",  x"21",  x"e1",  x"b7", -- 02E8
         x"cb",  x"4e",  x"20",  x"06",  x"ed",  x"53",  x"be",  x"b7", -- 02F0
         x"18",  x"04",  x"ed",  x"53",  x"c4",  x"b7",  x"c3",  x"8f", -- 02F8
         x"c3",  x"23",  x"46",  x"cd",  x"b1",  x"c3",  x"38",  x"32", -- 0300
         x"23",  x"23",  x"7e",  x"3d",  x"20",  x"0a",  x"3a",  x"e1", -- 0308
         x"b7",  x"cb",  x"97",  x"32",  x"e1",  x"b7",  x"18",  x"0b", -- 0310
         x"3d",  x"20",  x"1f",  x"3a",  x"e1",  x"b7",  x"cb",  x"d7", -- 0318
         x"32",  x"e1",  x"b7",  x"23",  x"23",  x"11",  x"06",  x"fa", -- 0320
         x"7e",  x"3d",  x"3d",  x"20",  x"0f",  x"ed",  x"53",  x"be", -- 0328
         x"b7",  x"11",  x"e1",  x"b7",  x"1a",  x"cb",  x"8f",  x"12", -- 0330
         x"18",  x"10",  x"18",  x"72",  x"3d",  x"20",  x"fb",  x"ed", -- 0338
         x"53",  x"c4",  x"b7",  x"11",  x"e1",  x"b7",  x"1a",  x"cb", -- 0340
         x"cf",  x"12",  x"3a",  x"81",  x"b7",  x"fe",  x"04",  x"23", -- 0348
         x"23",  x"38",  x"3c",  x"7e",  x"a7",  x"28",  x"1c",  x"3d", -- 0350
         x"28",  x"0a",  x"3d",  x"20",  x"51",  x"3a",  x"e1",  x"b7", -- 0358
         x"cb",  x"c7",  x"18",  x"05",  x"3a",  x"e1",  x"b7",  x"cb", -- 0360
         x"87",  x"32",  x"e1",  x"b7",  x"11",  x"e2",  x"f9",  x"ed", -- 0368
         x"53",  x"99",  x"b7",  x"3a",  x"81",  x"b7",  x"fe",  x"05", -- 0370
         x"20",  x"15",  x"23",  x"23",  x"7e",  x"cb",  x"27",  x"cb", -- 0378
         x"27",  x"cb",  x"27",  x"cb",  x"27",  x"4f",  x"3a",  x"e1", -- 0380
         x"b7",  x"e6",  x"0f",  x"b1",  x"32",  x"e1",  x"b7",  x"cd", -- 0388
         x"d4",  x"fa",  x"3e",  x"0c",  x"c5",  x"81",  x"06",  x"02", -- 0390
         x"4f",  x"2a",  x"e2",  x"b7",  x"f3",  x"ed",  x"b3",  x"c1", -- 0398
         x"3a",  x"e4",  x"b7",  x"3d",  x"3d",  x"47",  x"3e",  x"0a", -- 03A0
         x"81",  x"4f",  x"ed",  x"b3",  x"fb",  x"c9",  x"c3",  x"61", -- 03A8
         x"f3",  x"16",  x"3c",  x"0e",  x"80",  x"ed",  x"78",  x"fe", -- 03B0
         x"ee",  x"28",  x"09",  x"04",  x"04",  x"04",  x"04",  x"15", -- 03B8
         x"20",  x"f3",  x"37",  x"c9",  x"e5",  x"68",  x"3e",  x"02", -- 03C0
         x"16",  x"01",  x"cd",  x"04",  x"e4",  x"e1",  x"c9",  x"e5", -- 03C8
         x"d5",  x"3a",  x"e1",  x"b7",  x"cb",  x"47",  x"c2",  x"25", -- 03D0
         x"c4",  x"2a",  x"b9",  x"b7",  x"af",  x"b6",  x"20",  x"1a", -- 03D8
         x"11",  x"03",  x"fa",  x"3d",  x"3d",  x"28",  x"05",  x"21", -- 03E0
         x"a3",  x"fb",  x"18",  x"18",  x"21",  x"a2",  x"fb",  x"18", -- 03E8
         x"19",  x"ed",  x"53",  x"be",  x"b7",  x"21",  x"a2",  x"fb", -- 03F0
         x"18",  x"14",  x"3d",  x"11",  x"06",  x"fa",  x"21",  x"a0", -- 03F8
         x"fb",  x"3d",  x"28",  x"06",  x"ed",  x"53",  x"c4",  x"b7", -- 0400
         x"18",  x"04",  x"ed",  x"53",  x"be",  x"b7",  x"22",  x"b9", -- 0408
         x"b7",  x"d1",  x"e1",  x"c9",  x"1b",  x"5b",  x"31",  x"31", -- 0410
         x"61",  x"5b",  x"30",  x"31",  x"65",  x"1b",  x"5b",  x"37", -- 0418
         x"38",  x"71",  x"4b",  x"40",  x"02",  x"c5",  x"f5",  x"3a", -- 0420
         x"e1",  x"b7",  x"cb",  x"7f",  x"28",  x"2a",  x"2a",  x"cb", -- 0428
         x"b7",  x"06",  x"20",  x"0e",  x"28",  x"7e",  x"23",  x"a7", -- 0430
         x"20",  x"02",  x"3e",  x"20",  x"fe",  x"20",  x"30",  x"02", -- 0438
         x"3e",  x"20",  x"cd",  x"06",  x"fa",  x"0d",  x"20",  x"ed", -- 0440
         x"3e",  x"0d",  x"cd",  x"38",  x"fa",  x"3e",  x"0a",  x"cd", -- 0448
         x"38",  x"fa",  x"10",  x"df",  x"f1",  x"c3",  x"34",  x"f2", -- 0450
         x"e6",  x"f0",  x"28",  x"15",  x"fe",  x"10",  x"28",  x"5c", -- 0458
         x"fe",  x"20",  x"ca",  x"32",  x"c5",  x"fe",  x"30",  x"ca", -- 0460
         x"b7",  x"c5",  x"fe",  x"50",  x"ca",  x"fa",  x"c5",  x"18", -- 0468
         x"e3",  x"26",  x"00",  x"e5",  x"21",  x"16",  x"c6",  x"06", -- 0470
         x"0a",  x"cd",  x"0e",  x"c6",  x"e1",  x"cd",  x"8f",  x"c4", -- 0478
         x"30",  x"f1",  x"3e",  x"0d",  x"cd",  x"51",  x"fa",  x"3e", -- 0480
         x"0a",  x"cd",  x"51",  x"fa",  x"c3",  x"54",  x"c4",  x"2e", -- 0488
         x"00",  x"01",  x"08",  x"00",  x"e5",  x"11",  x"00",  x"b7", -- 0490
         x"cd",  x"4e",  x"e0",  x"ed",  x"b0",  x"0e",  x"08",  x"06", -- 0498
         x"08",  x"21",  x"00",  x"b7",  x"cb",  x"16",  x"17",  x"23", -- 04A0
         x"10",  x"fa",  x"cd",  x"51",  x"fa",  x"0d",  x"20",  x"ef", -- 04A8
         x"e1",  x"2c",  x"3e",  x"28",  x"bd",  x"20",  x"da",  x"7c", -- 04B0
         x"c6",  x"08",  x"67",  x"c9",  x"26",  x"00",  x"e5",  x"21", -- 04B8
         x"20",  x"c6",  x"06",  x"0a",  x"cd",  x"0e",  x"c6",  x"e1", -- 04C0
         x"2e",  x"00",  x"06",  x"04",  x"e5",  x"11",  x"00",  x"b7", -- 04C8
         x"cd",  x"4e",  x"e0",  x"7e",  x"12",  x"13",  x"12",  x"13", -- 04D0
         x"2c",  x"10",  x"f8",  x"0e",  x"08",  x"06",  x"08",  x"21", -- 04D8
         x"00",  x"b7",  x"cb",  x"16",  x"17",  x"23",  x"10",  x"fa", -- 04E0
         x"cd",  x"51",  x"fa",  x"cd",  x"51",  x"fa",  x"0d",  x"20", -- 04E8
         x"ec",  x"e1",  x"2c",  x"3e",  x"28",  x"bd",  x"20",  x"d2", -- 04F0
         x"7c",  x"c6",  x"04",  x"67",  x"30",  x"c0",  x"18",  x"82", -- 04F8
         x"e5",  x"c5",  x"cd",  x"4e",  x"e0",  x"06",  x"00",  x"ed", -- 0500
         x"b0",  x"c1",  x"e1",  x"c9",  x"e5",  x"c5",  x"2e",  x"80", -- 0508
         x"06",  x"00",  x"11",  x"00",  x"b7",  x"1a",  x"a5",  x"28", -- 0510
         x"01",  x"37",  x"cb",  x"10",  x"13",  x"3e",  x"06",  x"bb", -- 0518
         x"20",  x"f3",  x"a7",  x"cb",  x"10",  x"78",  x"cd",  x"51", -- 0520
         x"fa",  x"cb",  x"0d",  x"cb",  x"7d",  x"28",  x"e1",  x"c1", -- 0528
         x"e1",  x"c9",  x"21",  x"2a",  x"c6",  x"06",  x"0e",  x"cd", -- 0530
         x"0e",  x"c6",  x"06",  x"2a",  x"21",  x"00",  x"00",  x"11", -- 0538
         x"00",  x"b7",  x"0e",  x"06",  x"cd",  x"00",  x"c5",  x"cd", -- 0540
         x"0c",  x"c5",  x"2c",  x"3e",  x"28",  x"bd",  x"20",  x"ef", -- 0548
         x"3e",  x"06",  x"84",  x"67",  x"2e",  x"00",  x"e5",  x"c5", -- 0550
         x"21",  x"2a",  x"c6",  x"06",  x"0e",  x"cd",  x"0e",  x"c6", -- 0558
         x"c1",  x"e1",  x"05",  x"20",  x"da",  x"11",  x"00",  x"b7", -- 0560
         x"0e",  x"04",  x"cd",  x"00",  x"c5",  x"af",  x"12",  x"13", -- 0568
         x"12",  x"cd",  x"0c",  x"c5",  x"2c",  x"3e",  x"28",  x"bd", -- 0570
         x"20",  x"eb",  x"c3",  x"82",  x"c4",  x"e5",  x"11",  x"00", -- 0578
         x"b7",  x"cd",  x"4e",  x"e0",  x"7e",  x"12",  x"13",  x"12", -- 0580
         x"13",  x"2c",  x"0d",  x"20",  x"f7",  x"e1",  x"c9",  x"e5", -- 0588
         x"c5",  x"2e",  x"80",  x"06",  x"00",  x"11",  x"00",  x"b7", -- 0590
         x"1a",  x"a5",  x"28",  x"01",  x"37",  x"cb",  x"10",  x"13", -- 0598
         x"3e",  x"06",  x"bb",  x"20",  x"f3",  x"78",  x"17",  x"17", -- 05A0
         x"cd",  x"51",  x"fa",  x"cd",  x"51",  x"fa",  x"cb",  x"0d", -- 05A8
         x"cb",  x"7d",  x"28",  x"df",  x"c1",  x"e1",  x"c9",  x"21", -- 05B0
         x"38",  x"c6",  x"06",  x"0e",  x"cd",  x"0e",  x"c6",  x"06", -- 05B8
         x"55",  x"21",  x"00",  x"00",  x"0e",  x"03",  x"cd",  x"7d", -- 05C0
         x"c5",  x"cd",  x"8f",  x"c5",  x"2c",  x"3e",  x"28",  x"bd", -- 05C8
         x"20",  x"f2",  x"24",  x"24",  x"24",  x"2e",  x"00",  x"e5", -- 05D0
         x"c5",  x"21",  x"38",  x"c6",  x"06",  x"0e",  x"cd",  x"0e", -- 05D8
         x"c6",  x"c1",  x"e1",  x"10",  x"df",  x"0e",  x"01",  x"cd", -- 05E0
         x"7d",  x"c5",  x"af",  x"12",  x"13",  x"12",  x"cd",  x"8f", -- 05E8
         x"c5",  x"2c",  x"3e",  x"28",  x"bd",  x"20",  x"ee",  x"c3", -- 05F0
         x"82",  x"c4",  x"26",  x"00",  x"e5",  x"21",  x"46",  x"c6", -- 05F8
         x"06",  x"09",  x"cd",  x"0e",  x"c6",  x"e1",  x"cd",  x"8f", -- 0600
         x"c4",  x"30",  x"f1",  x"c3",  x"82",  x"c4",  x"7e",  x"23", -- 0608
         x"cd",  x"51",  x"fa",  x"10",  x"f9",  x"c9",  x"0d",  x"09", -- 0610
         x"1b",  x"4a",  x"18",  x"1b",  x"2a",  x"05",  x"40",  x"01", -- 0618
         x"0d",  x"09",  x"1b",  x"4a",  x"18",  x"1b",  x"2a",  x"05", -- 0620
         x"80",  x"02",  x"1b",  x"5b",  x"30",  x"31",  x"65",  x"1b", -- 0628
         x"5b",  x"31",  x"32",  x"60",  x"1b",  x"4b",  x"40",  x"01", -- 0630
         x"1b",  x"5b",  x"30",  x"31",  x"65",  x"1b",  x"5b",  x"31", -- 0638
         x"32",  x"60",  x"1b",  x"4b",  x"80",  x"02",  x"0d",  x"09", -- 0640
         x"1b",  x"4a",  x"18",  x"1b",  x"4b",  x"40",  x"01",  x"3a", -- 0648
         x"81",  x"b7",  x"fe",  x"03",  x"38",  x"29",  x"21",  x"82", -- 0650
         x"b7",  x"46",  x"cd",  x"b1",  x"c3",  x"da",  x"61",  x"f3", -- 0658
         x"23",  x"23",  x"3a",  x"e8",  x"b7",  x"cb",  x"46",  x"cb", -- 0660
         x"97",  x"20",  x"02",  x"cb",  x"d7",  x"47",  x"23",  x"23", -- 0668
         x"7e",  x"d6",  x"02",  x"cb",  x"88",  x"28",  x"02",  x"cb", -- 0670
         x"c8",  x"78",  x"32",  x"e8",  x"b7",  x"18",  x"06",  x"cd", -- 0678
         x"b1",  x"c3",  x"da",  x"61",  x"f3",  x"11",  x"78",  x"fa", -- 0680
         x"01",  x"98",  x"fa",  x"3a",  x"e8",  x"b7",  x"cb",  x"4f", -- 0688
         x"20",  x"0a",  x"ed",  x"53",  x"be",  x"b7",  x"ed",  x"43", -- 0690
         x"c1",  x"b7",  x"18",  x"08",  x"ed",  x"53",  x"c4",  x"b7", -- 0698
         x"ed",  x"43",  x"c7",  x"b7",  x"cd",  x"e1",  x"fa",  x"3e", -- 06A0
         x"0c",  x"c5",  x"81",  x"06",  x"02",  x"4f",  x"2a",  x"e5", -- 06A8
         x"b7",  x"f3",  x"ed",  x"b3",  x"c1",  x"3a",  x"e7",  x"b7", -- 06B0
         x"3d",  x"3d",  x"47",  x"3e",  x"0a",  x"81",  x"4f",  x"ed", -- 06B8
         x"b3",  x"fb",  x"c9",  x"21",  x"78",  x"fa",  x"22",  x"c4", -- 06C0
         x"b7",  x"0e",  x"0d",  x"21",  x"01",  x"c7",  x"06",  x"02", -- 06C8
         x"f3",  x"ed",  x"b3",  x"06",  x"0b",  x"0e",  x"0b",  x"18", -- 06D0
         x"e6",  x"21",  x"f0",  x"c6",  x"11",  x"01",  x"a8",  x"01", -- 06D8
         x"11",  x"00",  x"ed",  x"b0",  x"06",  x"08",  x"cd",  x"b1", -- 06E0
         x"c3",  x"d8",  x"3e",  x"01",  x"32",  x"00",  x"a8",  x"c9", -- 06E8
         x"47",  x"5b",  x"04",  x"04",  x"03",  x"20",  x"05",  x"6a", -- 06F0
         x"47",  x"2e",  x"18",  x"04",  x"44",  x"03",  x"e1",  x"05", -- 06F8
         x"6a",  x"47",  x"2e",  x"18",  x"02",  x"e2",  x"14",  x"44", -- 0700
         x"03",  x"e1",  x"05",  x"ea",  x"11",  x"18",  x"01",  x"81", -- 0708
         x"b7",  x"af",  x"02",  x"cd",  x"92",  x"f3",  x"d8",  x"7e", -- 0710
         x"b7",  x"c8",  x"23",  x"03",  x"7e",  x"02",  x"23",  x"03", -- 0718
         x"7e",  x"02",  x"2e",  x"81",  x"34",  x"7e",  x"c6",  x"f5", -- 0720
         x"30",  x"e9",  x"c9",  x"5a",  x"57",  x"d5",  x"c5",  x"cb", -- 0728
         x"5b",  x"28",  x"29",  x"dd",  x"cb",  x"07",  x"ce",  x"3e", -- 0730
         x"d5",  x"be",  x"d5",  x"11",  x"a0",  x"00",  x"20",  x"03", -- 0738
         x"11",  x"00",  x"05",  x"ed",  x"53",  x"d8",  x"b7",  x"11", -- 0740
         x"00",  x"b7",  x"01",  x"0b",  x"00",  x"ed",  x"b0",  x"eb", -- 0748
         x"d1",  x"72",  x"3e",  x"74",  x"cd",  x"9c",  x"c8",  x"c1", -- 0750
         x"d1",  x"cb",  x"9b",  x"c9",  x"2a",  x"da",  x"b7",  x"72", -- 0758
         x"cb",  x"73",  x"20",  x"23",  x"3a",  x"dc",  x"b7",  x"3d", -- 0760
         x"20",  x"ea",  x"dd",  x"cb",  x"07",  x"4e",  x"20",  x"08", -- 0768
         x"cd",  x"81",  x"c8",  x"cd",  x"95",  x"c8",  x"18",  x"df", -- 0770
         x"dd",  x"cb",  x"07",  x"8e",  x"cd",  x"1c",  x"e5",  x"cd", -- 0778
         x"88",  x"c8",  x"cd",  x"95",  x"c8",  x"18",  x"d0",  x"dd", -- 0780
         x"cb",  x"07",  x"4e",  x"28",  x"05",  x"cd",  x"1c",  x"e5", -- 0788
         x"18",  x"03",  x"cd",  x"81",  x"c8",  x"ed",  x"4b",  x"d8", -- 0790
         x"b7",  x"cd",  x"d9",  x"e4",  x"d5",  x"cd",  x"ff",  x"f5", -- 0798
         x"dd",  x"cb",  x"07",  x"ae",  x"d1",  x"18",  x"de",  x"5a", -- 07A0
         x"57",  x"d5",  x"c5",  x"cb",  x"73",  x"20",  x"ed",  x"cb", -- 07A8
         x"5b",  x"28",  x"66",  x"3e",  x"01",  x"dd",  x"77",  x"03", -- 07B0
         x"e5",  x"cd",  x"8e",  x"e5",  x"e1",  x"da",  x"71",  x"c8", -- 07B8
         x"dd",  x"7e",  x"02",  x"fe",  x"01",  x"c2",  x"71",  x"c8", -- 07C0
         x"dd",  x"cb",  x"07",  x"be",  x"dd",  x"34",  x"03",  x"11", -- 07C8
         x"00",  x"b7",  x"06",  x"0b",  x"1a",  x"fe",  x"d5",  x"20", -- 07D0
         x"04",  x"dd",  x"cb",  x"07",  x"ee",  x"c6",  x"29",  x"30", -- 07D8
         x"12",  x"1a",  x"d6",  x"04",  x"12",  x"13",  x"12",  x"13", -- 07E0
         x"12",  x"32",  x"5e",  x"03",  x"dd",  x"cb",  x"07",  x"f6", -- 07E8
         x"11",  x"00",  x"b7",  x"1a",  x"cd",  x"29",  x"e3",  x"be", -- 07F0
         x"28",  x"04",  x"dd",  x"cb",  x"07",  x"fe",  x"23",  x"13", -- 07F8
         x"10",  x"f1",  x"cd",  x"6b",  x"f3",  x"dd",  x"cb",  x"07", -- 0800
         x"7e",  x"c2",  x"7b",  x"f8",  x"eb",  x"3e",  x"75",  x"56", -- 0808
         x"cd",  x"9c",  x"c8",  x"7a",  x"c1",  x"d1",  x"cb",  x"9b", -- 0810
         x"c9",  x"2a",  x"da",  x"b7",  x"3a",  x"dc",  x"b7",  x"3d", -- 0818
         x"20",  x"ed",  x"cd",  x"91",  x"e5",  x"38",  x"39",  x"cd", -- 0820
         x"95",  x"c8",  x"3e",  x"ff",  x"dd",  x"be",  x"02",  x"28", -- 0828
         x"17",  x"dd",  x"7e",  x"03",  x"dd",  x"be",  x"02",  x"28", -- 0830
         x"0f",  x"3e",  x"2a",  x"cd",  x"29",  x"e3",  x"cd",  x"e8", -- 0838
         x"f1",  x"19",  x"00",  x"cd",  x"8e",  x"c8",  x"18",  x"da", -- 0840
         x"dd",  x"34",  x"03",  x"3d",  x"dd",  x"cb",  x"07",  x"6e", -- 0848
         x"20",  x"06",  x"cd",  x"e8",  x"f1",  x"3e",  x"19",  x"00", -- 0850
         x"cd",  x"95",  x"c8",  x"2a",  x"da",  x"b7",  x"18",  x"af", -- 0858
         x"cd",  x"ee",  x"f1",  x"09",  x"09",  x"09",  x"09",  x"3f", -- 0860
         x"00",  x"cd",  x"e8",  x"f1",  x"0d",  x"0a",  x"00",  x"18", -- 0868
         x"d2",  x"cd",  x"ee",  x"f1",  x"2a",  x"08",  x"00",  x"cd", -- 0870
         x"8e",  x"c8",  x"cd",  x"91",  x"e5",  x"e5",  x"c3",  x"bc", -- 0878
         x"c7",  x"ed",  x"4b",  x"d8",  x"b7",  x"cd",  x"2b",  x"e5", -- 0880
         x"cd",  x"e8",  x"f1",  x"3e",  x"19",  x"00",  x"cd",  x"de", -- 0888
         x"e3",  x"d0",  x"c3",  x"7b",  x"f8",  x"3e",  x"80",  x"21", -- 0890
         x"00",  x"b7",  x"18",  x"01",  x"23",  x"22",  x"da",  x"b7", -- 0898
         x"32",  x"dc",  x"b7",  x"c9",  x"00",  x"b9",  x"ca",  x"63", -- 08A0
         x"33",  x"c3",  x"79",  x"32",  x"04",  x"05",  x"ca",  x"87", -- 08A8
         x"33",  x"77",  x"2b",  x"04",  x"c3",  x"b2",  x"32",  x"05", -- 08B0
         x"ca",  x"b2",  x"32",  x"fa",  x"9a",  x"33",  x"c3",  x"b0", -- 08B8
         x"32",  x"04",  x"05",  x"c2",  x"b0",  x"32",  x"d1",  x"7b", -- 08C0
         x"95",  x"3d",  x"12",  x"c1",  x"eb",  x"2a",  x"2b",  x"3d", -- 08C8
         x"2b",  x"7e",  x"fe",  x"20",  x"cc",  x"30",  x"0b",  x"fe", -- 08D0
         x"09",  x"cc",  x"30",  x"0b",  x"eb",  x"c9",  x"04",  x"05", -- 08D8
         x"ca",  x"9a",  x"33",  x"cd",  x"df",  x"04",  x"c3",  x"9a", -- 08E0
         x"33",  x"f5",  x"e5",  x"21",  x"af",  x"3d",  x"cd",  x"87", -- 08E8
         x"0d",  x"d2",  x"d0",  x"33",  x"23",  x"36",  x"0d",  x"2b", -- 08F0
         x"eb",  x"e1",  x"f1",  x"c9",  x"e1",  x"f1",  x"12",  x"13", -- 08F8
         x"c9",  x"cd",  x"23",  x"31",  x"fe",  x"26",  x"ca",  x"d5", -- 0900
         x"33",  x"fe",  x"3a",  x"ca",  x"23",  x"31",  x"fe",  x"21", -- 0908
         x"d0",  x"fe",  x"0d",  x"c8",  x"f5",  x"cd",  x"08",  x"0c", -- 0910
         x"ca",  x"f5",  x"33",  x"cd",  x"0f",  x"05",  x"ca",  x"c1", -- 0918
         x"18",  x"f1",  x"c3",  x"23",  x"31",  x"21",  x"ff",  x"33", -- 0920
         x"c3",  x"6c",  x"0d",  x"3f",  x"53",  x"74",  x"61",  x"63", -- 0928
         x"6b",  x"20",  x"6f",  x"76",  x"65",  x"72",  x"66",  x"6c", -- 0930
         x"6f",  x"77",  x"2c",  x"20",  x"74",  x"72",  x"79",  x"20", -- 0938
         x"6d",  x"6f",  x"72",  x"65",  x"20",  x"50",  x"20",  x"73", -- 0940
         x"77",  x"69",  x"74",  x"63",  x"68",  x"65",  x"73",  x"0d", -- 0948
         x"0a",  x"00",  x"cd",  x"a9",  x"28",  x"3a",  x"f6",  x"3d", -- 0950
         x"fe",  x"20",  x"ca",  x"34",  x"34",  x"11",  x"00",  x"00", -- 0958
         x"eb",  x"22",  x"e2",  x"3f",  x"cd",  x"e3",  x"2f",  x"c1", -- 0960
         x"d1",  x"e1",  x"01",  x"48",  x"34",  x"c5",  x"d5",  x"3e", -- 0968
         x"0d",  x"c3",  x"56",  x"04",  x"c1",  x"01",  x"43",  x"34", -- 0970
         x"c5",  x"cd",  x"4f",  x"0b",  x"fe",  x"3a",  x"cc",  x"4f", -- 0978
         x"0b",  x"cd",  x"2d",  x"30",  x"ca",  x"69",  x"34",  x"11", -- 0980
         x"2d",  x"3d",  x"1a",  x"cd",  x"20",  x"3a",  x"13",  x"fe", -- 0988
         x"0d",  x"c2",  x"5e",  x"34",  x"c9",  x"af",  x"cd",  x"20", -- 0990
         x"3a",  x"cd",  x"83",  x"3a",  x"c1",  x"d1",  x"e1",  x"21", -- 0998
         x"cc",  x"02",  x"e5",  x"d5",  x"2a",  x"08",  x"40",  x"e5", -- 09A0
         x"e5",  x"2a",  x"e2",  x"3f",  x"e5",  x"21",  x"cc",  x"02", -- 09A8
         x"e5",  x"21",  x"8b",  x"34",  x"e5",  x"c5",  x"c9",  x"cd", -- 09B0
         x"de",  x"34",  x"c1",  x"e1",  x"d1",  x"cd",  x"87",  x"0d", -- 09B8
         x"c2",  x"ba",  x"34",  x"3a",  x"eb",  x"3f",  x"b7",  x"c2", -- 09C0
         x"a3",  x"34",  x"78",  x"b1",  x"c2",  x"ba",  x"34",  x"2a", -- 09C8
         x"dd",  x"3f",  x"e5",  x"cd",  x"79",  x"39",  x"e1",  x"cd", -- 09D0
         x"6f",  x"30",  x"af",  x"32",  x"eb",  x"3f",  x"d1",  x"d5", -- 09D8
         x"2a",  x"e4",  x"3f",  x"e5",  x"eb",  x"e9",  x"d5",  x"cd", -- 09E0
         x"57",  x"3a",  x"b7",  x"ca",  x"ed",  x"34",  x"11",  x"2d", -- 09E8
         x"3d",  x"cd",  x"6d",  x"3a",  x"cd",  x"bd",  x"33",  x"fe", -- 09F0
         x"0d",  x"c2",  x"c5",  x"34",  x"e5",  x"c5",  x"2a",  x"e6", -- 09F8
         x"3f",  x"e5",  x"2a",  x"e8",  x"3f",  x"e5",  x"2a",  x"e4", -- 0A00
         x"3f",  x"e9",  x"d1",  x"e1",  x"22",  x"e4",  x"3f",  x"e1", -- 0A08
         x"22",  x"e8",  x"3f",  x"e1",  x"22",  x"e6",  x"3f",  x"eb", -- 0A10
         x"e9",  x"0b",  x"62",  x"6b",  x"c3",  x"90",  x"34",  x"3a", -- 0A18
         x"df",  x"3f",  x"b7",  x"ca",  x"df",  x"04",  x"32",  x"eb", -- 0A20
         x"3f",  x"c1",  x"e1",  x"d1",  x"11",  x"10",  x"35",  x"d5", -- 0A28
         x"e5",  x"c5",  x"af",  x"32",  x"ea",  x"3f",  x"c3",  x"3a", -- 0A30
         x"0b",  x"c3",  x"bb",  x"04",  x"3a",  x"eb",  x"3f",  x"b7", -- 0A38
         x"ca",  x"6f",  x"35",  x"c1",  x"01",  x"de",  x"01",  x"c5", -- 0A40
         x"cd",  x"4f",  x"0b",  x"fe",  x"3a",  x"cc",  x"4f",  x"0b", -- 0A48
         x"cd",  x"0f",  x"05",  x"c0",  x"b7",  x"f0",  x"4f",  x"e6", -- 0A50
         x"08",  x"c2",  x"43",  x"35",  x"79",  x"e6",  x"10",  x"c2", -- 0A58
         x"4b",  x"35",  x"79",  x"e6",  x"20",  x"c2",  x"53",  x"35", -- 0A60
         x"79",  x"e6",  x"40",  x"c2",  x"60",  x"35",  x"c9",  x"3a", -- 0A68
         x"ea",  x"3f",  x"3d",  x"32",  x"ea",  x"3f",  x"c9",  x"3a", -- 0A70
         x"ea",  x"3f",  x"3c",  x"32",  x"ea",  x"3f",  x"c9",  x"3a", -- 0A78
         x"ea",  x"3f",  x"b7",  x"c0",  x"3a",  x"d8",  x"3c",  x"b7", -- 0A80
         x"c8",  x"c3",  x"cf",  x"28",  x"3a",  x"ea",  x"3f",  x"b7", -- 0A88
         x"c0",  x"23",  x"7e",  x"fe",  x"08",  x"c8",  x"3e",  x"ff", -- 0A90
         x"c3",  x"35",  x"29",  x"c1",  x"d1",  x"e1",  x"21",  x"cc", -- 0A98
         x"02",  x"e5",  x"d5",  x"c5",  x"c9",  x"b7",  x"f5",  x"cd", -- 0AA0
         x"e3",  x"2f",  x"22",  x"ec",  x"3f",  x"cd",  x"4e",  x"32", -- 0AA8
         x"4f",  x"3a",  x"f6",  x"3d",  x"fe",  x"20",  x"ca",  x"95", -- 0AB0
         x"35",  x"2a",  x"ec",  x"3f",  x"cd",  x"6f",  x"30",  x"f1", -- 0AB8
         x"c9",  x"79",  x"36",  x"00",  x"2b",  x"fe",  x"2c",  x"c4", -- 0AC0
         x"97",  x"04",  x"f1",  x"f5",  x"ca",  x"d1",  x"35",  x"cd", -- 0AC8
         x"23",  x"0b",  x"fe",  x"3c",  x"c4",  x"97",  x"04",  x"f1", -- 0AD0
         x"77",  x"e5",  x"f5",  x"0e",  x"00",  x"2b",  x"3a",  x"f6", -- 0AD8
         x"3d",  x"fe",  x"20",  x"c2",  x"2c",  x"36",  x"f1",  x"f5", -- 0AE0
         x"47",  x"ca",  x"df",  x"35",  x"cd",  x"71",  x"32",  x"0c", -- 0AE8
         x"fe",  x"0d",  x"ca",  x"29",  x"36",  x"fe",  x"3e",  x"ca", -- 0AF0
         x"2c",  x"36",  x"c3",  x"c0",  x"35",  x"cd",  x"1d",  x"0b", -- 0AF8
         x"d6",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0B98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0BA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0BA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0BB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0BB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0BC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0BC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0BD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0BD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0BE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0BE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0BF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0BF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0C98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0CA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0CA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0CB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0CB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0CC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0CC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0CD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0CD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0CE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0CE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0CF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0CF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0D98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0E98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0EA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0EA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0EB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0EB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0EC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0EC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0ED0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0ED8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0EE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0EE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0EF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0EF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0F98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FF0
         x"ff",  x"ff",  x"5c",  x"98",  x"01",  x"1c",  x"d5",  x"79"  -- 0FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
