library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity caos47_c is
    generic(
        ADDR_WIDTH   : integer := 13
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end caos47_c;

architecture rtl of caos47_c is
    type rom8192x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom8192x8 := (
         x"bf",  x"f4",  x"00",  x"00",  x"00",  x"28",  x"20",  x"00", -- 0000
         x"00",  x"00",  x"39",  x"69",  x"e2",  x"00",  x"ee",  x"00", -- 0008
         x"fe",  x"00",  x"ee",  x"00",  x"fe",  x"c4",  x"01",  x"00", -- 0010
         x"aa",  x"8f",  x"fc",  x"d3",  x"88",  x"c3",  x"12",  x"f0", -- 0018
         x"05",  x"f0",  x"0e",  x"f0",  x"c3",  x"bf",  x"f4",  x"c3", -- 0020
         x"bf",  x"f4",  x"c3",  x"bf",  x"f4",  x"c3",  x"bf",  x"f4", -- 0028
         x"82",  x"dc",  x"00",  x"b2",  x"47",  x"0c",  x"b5",  x"ed", -- 0030
         x"0e",  x"05",  x"00",  x"01",  x"a8",  x"08",  x"09",  x"a8", -- 0038
         x"09",  x"ee",  x"c3",  x"bf",  x"f4",  x"25",  x"ff",  x"d8", -- 0040
         x"ef",  x"94",  x"aa",  x"03",  x"01",  x"00",  x"03",  x"03", -- 0048
         x"00",  x"f3",  x"31",  x"00",  x"c0",  x"01",  x"00",  x"60", -- 0050
         x"61",  x"69",  x"e5",  x"0d",  x"20",  x"fc",  x"10",  x"fa", -- 0058
         x"31",  x"c4",  x"01",  x"0e",  x"80",  x"ed",  x"69",  x"10", -- 0060
         x"fc",  x"cd",  x"91",  x"c0",  x"21",  x"59",  x"d9",  x"11", -- 0068
         x"94",  x"aa",  x"01",  x"0c",  x"00",  x"ed",  x"b0",  x"af", -- 0070
         x"32",  x"9b",  x"b7",  x"cd",  x"e7",  x"c5",  x"3c",  x"fe", -- 0078
         x"0a",  x"38",  x"f5",  x"cd",  x"61",  x"f9",  x"3e",  x"0c", -- 0080
         x"cd",  x"8c",  x"e0",  x"cd",  x"57",  x"f9",  x"c3",  x"70", -- 0088
         x"f1",  x"f3",  x"ed",  x"5e",  x"21",  x"25",  x"d9",  x"cd", -- 0090
         x"58",  x"f5",  x"dd",  x"21",  x"f0",  x"01",  x"dd",  x"36", -- 0098
         x"01",  x"28",  x"dd",  x"36",  x"04",  x"e3",  x"dd",  x"36", -- 00A0
         x"08",  x"80",  x"11",  x"99",  x"b7",  x"21",  x"00",  x"c0", -- 00A8
         x"01",  x"34",  x"00",  x"ed",  x"b0",  x"1e",  x"db",  x"0e", -- 00B0
         x"17",  x"ed",  x"b0",  x"11",  x"00",  x"b8",  x"3a",  x"04", -- 00B8
         x"b8",  x"e6",  x"04",  x"0e",  x"06",  x"ed",  x"b0",  x"21", -- 00C0
         x"04",  x"b8",  x"b6",  x"77",  x"11",  x"00",  x"aa",  x"21", -- 00C8
         x"51",  x"d8",  x"01",  x"94",  x"00",  x"ed",  x"b0",  x"11", -- 00D0
         x"00",  x"a9",  x"3e",  x"08",  x"21",  x"e5",  x"d8",  x"01", -- 00D8
         x"20",  x"00",  x"ed",  x"b0",  x"3d",  x"20",  x"f5",  x"32", -- 00E0
         x"00",  x"a9",  x"11",  x"20",  x"a9",  x"01",  x"80",  x"fc", -- 00E8
         x"ed",  x"78",  x"fe",  x"a7",  x"20",  x"15",  x"3e",  x"04", -- 00F0
         x"32",  x"fc",  x"b8",  x"ed",  x"79",  x"01",  x"f3",  x"b3", -- 00F8
         x"ed",  x"78",  x"fe",  x"05",  x"20",  x"05",  x"01",  x"20", -- 0100
         x"00",  x"ed",  x"b0",  x"06",  x"08",  x"0e",  x"80",  x"ed", -- 0108
         x"78",  x"fe",  x"fd",  x"28",  x"09",  x"fe",  x"f9",  x"28", -- 0110
         x"05",  x"04",  x"20",  x"f3",  x"18",  x"34",  x"c5",  x"68", -- 0118
         x"cd",  x"62",  x"c3",  x"7e",  x"23",  x"be",  x"20",  x"1a", -- 0120
         x"fe",  x"46",  x"20",  x"16",  x"23",  x"7b",  x"07",  x"07", -- 0128
         x"07",  x"12",  x"13",  x"e3",  x"7c",  x"12",  x"13",  x"e3", -- 0130
         x"01",  x"1e",  x"00",  x"ed",  x"b0",  x"21",  x"e3",  x"ff", -- 0138
         x"19",  x"7e",  x"c1",  x"c5",  x"d5",  x"cc",  x"6d",  x"ed", -- 0140
         x"cd",  x"7b",  x"c3",  x"d1",  x"c1",  x"7a",  x"fe",  x"aa", -- 0148
         x"20",  x"c7",  x"3a",  x"20",  x"a9",  x"fe",  x"01",  x"cc", -- 0150
         x"f2",  x"d5",  x"3e",  x"01",  x"21",  x"65",  x"d9",  x"f3", -- 0158
         x"32",  x"d7",  x"b7",  x"ed",  x"47",  x"ed",  x"5e",  x"1e", -- 0160
         x"e0",  x"57",  x"01",  x"10",  x"00",  x"ed",  x"b0",  x"dd", -- 0168
         x"66",  x"01",  x"dd",  x"6e",  x"04",  x"dd",  x"7e",  x"08", -- 0170
         x"d5",  x"dd",  x"e1",  x"dd",  x"77",  x"08",  x"dd",  x"74", -- 0178
         x"01",  x"dd",  x"75",  x"04",  x"dd",  x"36",  x"0e",  x"0f", -- 0180
         x"dd",  x"36",  x"0f",  x"fc",  x"dd",  x"36",  x"09",  x"7f", -- 0188
         x"21",  x"3f",  x"d9",  x"cd",  x"58",  x"f5",  x"21",  x"9d", -- 0190
         x"ed",  x"cd",  x"58",  x"f5",  x"cd",  x"46",  x"f5",  x"fb", -- 0198
         x"c9",  x"2e",  x"ff",  x"cd",  x"cf",  x"f0",  x"2d",  x"2d", -- 01A0
         x"20",  x"2d",  x"2d",  x"20",  x"2d",  x"2d",  x"20",  x"43", -- 01A8
         x"41",  x"4f",  x"53",  x"45",  x"00",  x"db",  x"88",  x"e6", -- 01B0
         x"01",  x"18",  x"3b",  x"3e",  x"01",  x"cd",  x"9c",  x"c3", -- 01B8
         x"cd",  x"4e",  x"d3",  x"7d",  x"a7",  x"20",  x"12",  x"cd", -- 01C0
         x"cf",  x"f0",  x"52",  x"41",  x"4d",  x"30",  x"00",  x"db", -- 01C8
         x"88",  x"e6",  x"0f",  x"fe",  x"08",  x"cb",  x"4f",  x"18", -- 01D0
         x"1d",  x"3d",  x"20",  x"1c",  x"cd",  x"cf",  x"f0",  x"42", -- 01D8
         x"49",  x"4c",  x"44",  x"20",  x"00",  x"dd",  x"7e",  x"01", -- 01E0
         x"e6",  x"04",  x"0f",  x"0f",  x"c6",  x"30",  x"cd",  x"d5", -- 01E8
         x"f3",  x"3a",  x"01",  x"b8",  x"e6",  x"01",  x"18",  x"72", -- 01F0
         x"3d",  x"20",  x"1c",  x"cd",  x"cf",  x"f0",  x"55",  x"53", -- 01F8
         x"45",  x"52",  x"20",  x"00",  x"dd",  x"7e",  x"04",  x"07", -- 0200
         x"07",  x"07",  x"e6",  x"03",  x"ee",  x"33",  x"cd",  x"d5", -- 0208
         x"f3",  x"db",  x"88",  x"e6",  x"80",  x"18",  x"53",  x"3d", -- 0210
         x"20",  x"1e",  x"cd",  x"cf",  x"f0",  x"52",  x"41",  x"4d", -- 0218
         x"38",  x"20",  x"00",  x"dd",  x"7e",  x"01",  x"0f",  x"0f", -- 0220
         x"0f",  x"0f",  x"d6",  x"02",  x"cd",  x"cd",  x"f3",  x"db", -- 0228
         x"89",  x"cb",  x"6f",  x"07",  x"07",  x"3f",  x"18",  x"32", -- 0230
         x"3d",  x"20",  x"21",  x"cd",  x"cf",  x"f0",  x"52",  x"41", -- 0238
         x"4d",  x"34",  x"00",  x"cd",  x"bc",  x"f3",  x"3a",  x"04", -- 0240
         x"b8",  x"0f",  x"0f",  x"e6",  x"01",  x"c6",  x"30",  x"cd", -- 0248
         x"d5",  x"f3",  x"dd",  x"7e",  x"04",  x"cb",  x"47",  x"0f", -- 0250
         x"0f",  x"3f",  x"18",  x"0e",  x"cd",  x"cf",  x"f0",  x"43", -- 0258
         x"41",  x"4f",  x"53",  x"43",  x"00",  x"3a",  x"05",  x"b8", -- 0260
         x"e6",  x"01",  x"cd",  x"2d",  x"d3",  x"2c",  x"3e",  x"06", -- 0268
         x"bd",  x"c2",  x"bb",  x"c1",  x"c9",  x"af",  x"d3",  x"91", -- 0270
         x"db",  x"91",  x"a7",  x"20",  x"16",  x"cd",  x"cf",  x"f0", -- 0278
         x"2d",  x"2d",  x"20",  x"2d",  x"2d",  x"20",  x"2d",  x"2d", -- 0280
         x"20",  x"4a",  x"4f",  x"59",  x"2f",  x"43",  x"45",  x"4e", -- 0288
         x"0d",  x"0a",  x"00",  x"2e",  x"07",  x"e5",  x"3e",  x"01", -- 0290
         x"cd",  x"9c",  x"c3",  x"7c",  x"3c",  x"28",  x"36",  x"cd", -- 0298
         x"4e",  x"d3",  x"4c",  x"7c",  x"fe",  x"f3",  x"28",  x"32", -- 02A0
         x"fe",  x"fb",  x"28",  x"45",  x"fe",  x"fd",  x"ca",  x"15", -- 02A8
         x"c3",  x"21",  x"ae",  x"cf",  x"fe",  x"c0",  x"38",  x"04", -- 02B0
         x"fe",  x"d8",  x"38",  x"13",  x"21",  x"72",  x"ce",  x"7e", -- 02B8
         x"23",  x"fe",  x"ff",  x"28",  x"0a",  x"b9",  x"28",  x"07", -- 02C0
         x"7e",  x"23",  x"a7",  x"20",  x"fb",  x"18",  x"f0",  x"cd", -- 02C8
         x"06",  x"f9",  x"cd",  x"db",  x"f4",  x"e1",  x"2c",  x"20", -- 02D0
         x"bc",  x"c9",  x"cd",  x"62",  x"c3",  x"7e",  x"34",  x"be", -- 02D8
         x"77",  x"21",  x"c4",  x"cf",  x"28",  x"03",  x"21",  x"bb", -- 02E0
         x"cf",  x"cd",  x"06",  x"f9",  x"cd",  x"7b",  x"c3",  x"18", -- 02E8
         x"e1",  x"cd",  x"62",  x"c3",  x"11",  x"ad",  x"cf",  x"01", -- 02F0
         x"00",  x"20",  x"cd",  x"57",  x"f3",  x"38",  x"05",  x"21", -- 02F8
         x"a5",  x"cf",  x"18",  x"07",  x"2b",  x"7e",  x"fe",  x"7f", -- 0300
         x"20",  x"fa",  x"23",  x"7e",  x"fe",  x"20",  x"38",  x"dc", -- 0308
         x"cd",  x"d5",  x"f3",  x"18",  x"f5",  x"26",  x"b8",  x"7e", -- 0310
         x"cb",  x"d7",  x"45",  x"0e",  x"80",  x"ed",  x"79",  x"21", -- 0318
         x"b3",  x"cf",  x"db",  x"28",  x"3c",  x"20",  x"08",  x"db", -- 0320
         x"29",  x"3c",  x"20",  x"03",  x"21",  x"b7",  x"cf",  x"18", -- 0328
         x"b8",  x"53",  x"fe",  x"01",  x"f5",  x"28",  x"0d",  x"2d", -- 0330
         x"20",  x"09",  x"2c",  x"26",  x"b8",  x"5e",  x"72",  x"26", -- 0338
         x"ff",  x"18",  x"05",  x"2c",  x"cd",  x"9c",  x"c3",  x"5f", -- 0340
         x"cd",  x"b8",  x"f3",  x"7c",  x"cd",  x"b9",  x"f3",  x"7b", -- 0348
         x"cd",  x"c4",  x"f3",  x"f1",  x"28",  x"09",  x"3e",  x"09", -- 0350
         x"cd",  x"b5",  x"f7",  x"7a",  x"cd",  x"c4",  x"f3",  x"c3", -- 0358
         x"db",  x"f4",  x"01",  x"80",  x"08",  x"af",  x"ed",  x"79", -- 0360
         x"04",  x"7d",  x"b8",  x"20",  x"f8",  x"3e",  x"41",  x"ed", -- 0368
         x"79",  x"dd",  x"cb",  x"04",  x"87",  x"d3",  x"86",  x"21", -- 0370
         x"00",  x"40",  x"c9",  x"21",  x"04",  x"b8",  x"56",  x"e5", -- 0378
         x"3e",  x"02",  x"cd",  x"9c",  x"c3",  x"e1",  x"2c",  x"20", -- 0380
         x"f5",  x"c9",  x"0e",  x"80",  x"ed",  x"78",  x"fe",  x"ee", -- 0388
         x"28",  x"05",  x"04",  x"20",  x"f7",  x"37",  x"c9",  x"68", -- 0390
         x"3e",  x"02",  x"16",  x"01",  x"26",  x"b8",  x"0e",  x"80", -- 0398
         x"45",  x"fe",  x"02",  x"7e",  x"30",  x"04",  x"56",  x"ed", -- 03A0
         x"60",  x"c9",  x"f5",  x"72",  x"67",  x"7d",  x"fe",  x"06", -- 03A8
         x"38",  x"05",  x"ed",  x"51",  x"f1",  x"18",  x"f0",  x"04", -- 03B0
         x"f3",  x"db",  x"88",  x"10",  x"0d",  x"e6",  x"f5",  x"67", -- 03B8
         x"7a",  x"0f",  x"e6",  x"81",  x"17",  x"17",  x"07",  x"b4", -- 03C0
         x"18",  x"25",  x"10",  x"0a",  x"e6",  x"fb",  x"cb",  x"42", -- 03C8
         x"28",  x"1d",  x"f6",  x"04",  x"18",  x"19",  x"10",  x"1b", -- 03D0
         x"7a",  x"2f",  x"07",  x"e6",  x"60",  x"67",  x"dd",  x"7e", -- 03D8
         x"04",  x"e6",  x"9f",  x"b4",  x"dd",  x"77",  x"04",  x"d3", -- 03E0
         x"86",  x"7a",  x"0f",  x"db",  x"88",  x"17",  x"0f",  x"d3", -- 03E8
         x"88",  x"18",  x"23",  x"10",  x"26",  x"3e",  x"03",  x"a2", -- 03F0
         x"0f",  x"0f",  x"0f",  x"67",  x"db",  x"89",  x"e6",  x"9f", -- 03F8
         x"b4",  x"d3",  x"89",  x"7a",  x"07",  x"07",  x"c6",  x"20", -- 0400
         x"e6",  x"f0",  x"67",  x"dd",  x"7e",  x"01",  x"e6",  x"0f", -- 0408
         x"b4",  x"d3",  x"84",  x"dd",  x"77",  x"01",  x"fb",  x"f1", -- 0410
         x"26",  x"ff",  x"c9",  x"10",  x"f9",  x"7a",  x"ac",  x"e6", -- 0418
         x"04",  x"28",  x"3f",  x"dd",  x"7e",  x"04",  x"f6",  x"03", -- 0420
         x"d3",  x"86",  x"d5",  x"e5",  x"db",  x"88",  x"f5",  x"cb", -- 0428
         x"87",  x"d3",  x"88",  x"dd",  x"7e",  x"01",  x"f5",  x"e6", -- 0430
         x"f9",  x"2e",  x"03",  x"01",  x"00",  x"10",  x"11",  x"00", -- 0438
         x"40",  x"c6",  x"02",  x"d3",  x"84",  x"67",  x"e5",  x"21", -- 0440
         x"00",  x"a8",  x"1a",  x"ed",  x"a0",  x"2b",  x"77",  x"23", -- 0448
         x"ea",  x"4a",  x"c4",  x"e1",  x"7c",  x"06",  x"18",  x"2d", -- 0450
         x"20",  x"e7",  x"f1",  x"d3",  x"84",  x"f1",  x"d3",  x"88", -- 0458
         x"e1",  x"d1",  x"dd",  x"7e",  x"04",  x"aa",  x"e6",  x"fc", -- 0460
         x"aa",  x"dd",  x"77",  x"04",  x"d3",  x"86",  x"18",  x"a6", -- 0468
         x"21",  x"00",  x"b9",  x"a7",  x"20",  x"07",  x"06",  x"9c", -- 0470
         x"77",  x"2c",  x"10",  x"fc",  x"c9",  x"fe",  x"10",  x"d0", -- 0478
         x"47",  x"f6",  x"f0",  x"4f",  x"7e",  x"2c",  x"c8",  x"a7", -- 0480
         x"20",  x"fa",  x"10",  x"f8",  x"7d",  x"fe",  x"9c",  x"d0", -- 0488
         x"ed",  x"5b",  x"a0",  x"b7",  x"cd",  x"4d",  x"c5",  x"cd", -- 0490
         x"f0",  x"f3",  x"fe",  x"13",  x"20",  x"03",  x"04",  x"18", -- 0498
         x"f6",  x"cb",  x"40",  x"28",  x"0d",  x"fe",  x"03",  x"28", -- 04A0
         x"70",  x"fe",  x"0d",  x"28",  x"0a",  x"cd",  x"d5",  x"f3", -- 04A8
         x"18",  x"e5",  x"cd",  x"b5",  x"f7",  x"18",  x"e0",  x"e5", -- 04B0
         x"cd",  x"68",  x"e0",  x"eb",  x"cd",  x"eb",  x"f4",  x"e1", -- 04B8
         x"38",  x"06",  x"3a",  x"97",  x"b7",  x"b9",  x"28",  x"06", -- 04C0
         x"cd",  x"db",  x"f4",  x"c3",  x"d1",  x"f4",  x"13",  x"13", -- 04C8
         x"06",  x"9b",  x"2f",  x"a7",  x"28",  x"21",  x"3c",  x"47", -- 04D0
         x"4d",  x"7e",  x"2c",  x"28",  x"eb",  x"a7",  x"20",  x"f9", -- 04D8
         x"10",  x"f7",  x"2d",  x"7d",  x"fe",  x"9c",  x"30",  x"e0", -- 04E0
         x"44",  x"c5",  x"91",  x"4f",  x"06",  x"00",  x"d5",  x"11", -- 04E8
         x"9b",  x"b9",  x"ed",  x"b8",  x"43",  x"d1",  x"e1",  x"4f", -- 04F0
         x"2d",  x"7e",  x"a7",  x"20",  x"fb",  x"2c",  x"1a",  x"13", -- 04F8
         x"77",  x"b7",  x"28",  x"08",  x"78",  x"95",  x"20",  x"f5", -- 0500
         x"36",  x"00",  x"18",  x"bc",  x"79",  x"a7",  x"28",  x"09", -- 0508
         x"04",  x"2c",  x"5d",  x"54",  x"68",  x"06",  x"00",  x"ed", -- 0510
         x"b0",  x"c3",  x"db",  x"f4",  x"21",  x"01",  x"b9",  x"01", -- 0518
         x"f1",  x"00",  x"7e",  x"a7",  x"28",  x"07",  x"cd",  x"4d", -- 0520
         x"c5",  x"cd",  x"db",  x"f4",  x"04",  x"2c",  x"7d",  x"fe", -- 0528
         x"9c",  x"30",  x"03",  x"0c",  x"20",  x"ec",  x"04",  x"05", -- 0530
         x"c0",  x"cd",  x"cf",  x"f0",  x"46",  x"2d",  x"54",  x"61", -- 0538
         x"73",  x"74",  x"65",  x"6e",  x"20",  x"6c",  x"65",  x"65", -- 0540
         x"72",  x"0d",  x"0a",  x"00",  x"c9",  x"3e",  x"02",  x"cd", -- 0548
         x"d5",  x"f3",  x"79",  x"cd",  x"cc",  x"f0",  x"20",  x"3a", -- 0550
         x"00",  x"7e",  x"b7",  x"c8",  x"cd",  x"b5",  x"f7",  x"23", -- 0558
         x"7d",  x"fe",  x"9c",  x"d0",  x"18",  x"f3",  x"a7",  x"20", -- 0560
         x"17",  x"3a",  x"a3",  x"b7",  x"6f",  x"0f",  x"0f",  x"0f", -- 0568
         x"e6",  x"1f",  x"cd",  x"b9",  x"f3",  x"7d",  x"e6",  x"07", -- 0570
         x"cd",  x"c4",  x"f3",  x"cd",  x"db",  x"f4",  x"18",  x"18", -- 0578
         x"3e",  x"1f",  x"a5",  x"17",  x"17",  x"17",  x"6f",  x"3a", -- 0580
         x"81",  x"b7",  x"fe",  x"02",  x"7b",  x"30",  x"03",  x"3a", -- 0588
         x"a3",  x"b7",  x"e6",  x"07",  x"b5",  x"32",  x"a3",  x"b7", -- 0590
         x"c3",  x"9c",  x"fb",  x"a7",  x"28",  x"20",  x"3d",  x"7d", -- 0598
         x"28",  x"28",  x"65",  x"69",  x"53",  x"3a",  x"88",  x"b7", -- 05A0
         x"5f",  x"3a",  x"81",  x"b7",  x"fe",  x"04",  x"38",  x"0b", -- 05A8
         x"3e",  x"00",  x"28",  x"03",  x"3a",  x"8a",  x"b7",  x"cd", -- 05B0
         x"fa",  x"c5",  x"d0",  x"c3",  x"d1",  x"f4",  x"11",  x"9b", -- 05B8
         x"b7",  x"21",  x"02",  x"c0",  x"01",  x"0b",  x"00",  x"ed", -- 05C0
         x"b0",  x"c9",  x"cd",  x"e7",  x"c5",  x"32",  x"9b",  x"b7", -- 05C8
         x"cd",  x"da",  x"c5",  x"d8",  x"eb",  x"11",  x"9c",  x"b7", -- 05D0
         x"18",  x"1a",  x"c6",  x"f6",  x"d8",  x"87",  x"5f",  x"87", -- 05D8
         x"87",  x"83",  x"5f",  x"16",  x"b9",  x"a7",  x"c9",  x"f5", -- 05E0
         x"3a",  x"9b",  x"b7",  x"cd",  x"da",  x"c5",  x"38",  x"3d", -- 05E8
         x"f1",  x"21",  x"9c",  x"b7",  x"01",  x"0a",  x"00",  x"ed", -- 05F0
         x"b0",  x"c9",  x"f5",  x"fe",  x"0a",  x"30",  x"2e",  x"7a", -- 05F8
         x"a7",  x"28",  x"2a",  x"84",  x"38",  x"27",  x"fe",  x"21", -- 0600
         x"30",  x"23",  x"7b",  x"a7",  x"28",  x"1f",  x"85",  x"38", -- 0608
         x"1c",  x"fe",  x"29",  x"30",  x"18",  x"f1",  x"d5",  x"e5", -- 0610
         x"cd",  x"e7",  x"c5",  x"e1",  x"d1",  x"22",  x"9c",  x"b7", -- 0618
         x"ed",  x"53",  x"9e",  x"b7",  x"ed",  x"43",  x"a0",  x"b7", -- 0620
         x"32",  x"9b",  x"b7",  x"a7",  x"c9",  x"f1",  x"37",  x"c9", -- 0628
         x"ed",  x"5b",  x"84",  x"b7",  x"2a",  x"88",  x"b7",  x"d9", -- 0630
         x"ed",  x"5b",  x"82",  x"b7",  x"d5",  x"2a",  x"86",  x"b7", -- 0638
         x"3e",  x"08",  x"b7",  x"ed",  x"52",  x"30",  x"06",  x"19", -- 0640
         x"eb",  x"f6",  x"01",  x"ed",  x"52",  x"d9",  x"d5",  x"ed", -- 0648
         x"52",  x"30",  x"06",  x"19",  x"eb",  x"f6",  x"02",  x"ed", -- 0650
         x"52",  x"e5",  x"d9",  x"c1",  x"e5",  x"ed",  x"42",  x"e1", -- 0658
         x"c5",  x"30",  x"05",  x"e3",  x"cb",  x"9f",  x"cb",  x"d7", -- 0660
         x"e5",  x"44",  x"4d",  x"d9",  x"c1",  x"d1",  x"60",  x"69", -- 0668
         x"cb",  x"3c",  x"cb",  x"1d",  x"d9",  x"d1",  x"e1",  x"f5", -- 0670
         x"08",  x"f1",  x"e5",  x"21",  x"ed",  x"b7",  x"cb",  x"06", -- 0678
         x"e1",  x"dc",  x"1e",  x"c7",  x"d9",  x"a7",  x"ed",  x"52", -- 0680
         x"30",  x"01",  x"09",  x"d9",  x"30",  x"02",  x"f6",  x"0c", -- 0688
         x"cb",  x"5f",  x"28",  x"07",  x"23",  x"cb",  x"47",  x"28", -- 0690
         x"02",  x"2b",  x"2b",  x"cb",  x"57",  x"28",  x"07",  x"13", -- 0698
         x"cb",  x"4f",  x"28",  x"02",  x"1b",  x"1b",  x"78",  x"b1", -- 06A0
         x"c8",  x"0b",  x"08",  x"18",  x"ca",  x"3a",  x"86",  x"b7", -- 06A8
         x"4f",  x"51",  x"cd",  x"db",  x"d2",  x"60",  x"6f",  x"54", -- 06B0
         x"5d",  x"79",  x"06",  x"00",  x"cb",  x"21",  x"cb",  x"10", -- 06B8
         x"0b",  x"c5",  x"01",  x"01",  x"00",  x"d9",  x"4f",  x"06", -- 06C0
         x"00",  x"e5",  x"21",  x"ed",  x"b7",  x"cb",  x"06",  x"e1", -- 06C8
         x"30",  x"06",  x"cd",  x"f8",  x"c6",  x"cd",  x"f8",  x"c6", -- 06D0
         x"d9",  x"a7",  x"ed",  x"42",  x"03",  x"03",  x"ed",  x"52", -- 06D8
         x"19",  x"d9",  x"30",  x"0c",  x"d9",  x"e3",  x"eb",  x"a7", -- 06E0
         x"ed",  x"52",  x"1b",  x"1b",  x"eb",  x"e3",  x"d9",  x"0d", -- 06E8
         x"04",  x"79",  x"b8",  x"30",  x"d4",  x"f1",  x"b7",  x"c9", -- 06F0
         x"78",  x"41",  x"4f",  x"af",  x"57",  x"2a",  x"84",  x"b7", -- 06F8
         x"e5",  x"59",  x"19",  x"cd",  x"0c",  x"c7",  x"af",  x"57", -- 0700
         x"e1",  x"59",  x"ed",  x"52",  x"e5",  x"2a",  x"82",  x"b7", -- 0708
         x"58",  x"a7",  x"ed",  x"52",  x"d1",  x"cd",  x"1e",  x"c7", -- 0710
         x"d5",  x"57",  x"58",  x"19",  x"19",  x"d1",  x"e5",  x"d5", -- 0718
         x"c5",  x"f5",  x"cd",  x"cd",  x"c7",  x"d4",  x"2b",  x"c7", -- 0720
         x"c3",  x"97",  x"e0",  x"dd",  x"cb",  x"01",  x"5e",  x"28", -- 0728
         x"29",  x"cb",  x"4a",  x"20",  x"21",  x"cb",  x"42",  x"20", -- 0730
         x"03",  x"b6",  x"18",  x"03",  x"ae",  x"cb",  x"82",  x"77", -- 0738
         x"cb",  x"52",  x"c0",  x"dd",  x"7e",  x"01",  x"5f",  x"ee", -- 0740
         x"02",  x"f3",  x"d3",  x"84",  x"7e",  x"e6",  x"07",  x"b2", -- 0748
         x"77",  x"7b",  x"d3",  x"84",  x"fb",  x"c9",  x"2f",  x"a6", -- 0750
         x"77",  x"c9",  x"47",  x"b6",  x"cb",  x"5a",  x"20",  x"01", -- 0758
         x"a8",  x"77",  x"dd",  x"7e",  x"01",  x"5f",  x"ee",  x"02", -- 0760
         x"f3",  x"d3",  x"84",  x"78",  x"b6",  x"cb",  x"62",  x"20", -- 0768
         x"df",  x"a8",  x"18",  x"dc",  x"e5",  x"d5",  x"c5",  x"cd", -- 0770
         x"c4",  x"c7",  x"d4",  x"2b",  x"c7",  x"18",  x"42",  x"e5", -- 0778
         x"d5",  x"c5",  x"cd",  x"c4",  x"c7",  x"38",  x"3a",  x"dd", -- 0780
         x"cb",  x"01",  x"5e",  x"20",  x"1e",  x"16",  x"00",  x"47", -- 0788
         x"7e",  x"a0",  x"28",  x"02",  x"cb",  x"c2",  x"dd",  x"7e", -- 0790
         x"01",  x"5f",  x"ee",  x"02",  x"f3",  x"d3",  x"84",  x"7e", -- 0798
         x"a0",  x"cd",  x"51",  x"c7",  x"28",  x"02",  x"cb",  x"ca", -- 07A0
         x"04",  x"18",  x"15",  x"47",  x"4e",  x"2f",  x"a1",  x"77", -- 07A8
         x"dd",  x"7e",  x"01",  x"5f",  x"ee",  x"02",  x"f3",  x"d3", -- 07B0
         x"84",  x"56",  x"7b",  x"d3",  x"84",  x"fb",  x"78",  x"a1", -- 07B8
         x"7a",  x"c3",  x"ec",  x"f3",  x"2a",  x"d3",  x"b7",  x"ed", -- 07C0
         x"5b",  x"d5",  x"b7",  x"16",  x"00",  x"c5",  x"01",  x"f8", -- 07C8
         x"fd",  x"7d",  x"e6",  x"07",  x"81",  x"4f",  x"7d",  x"cb", -- 07D0
         x"3c",  x"1f",  x"cb",  x"3c",  x"1f",  x"cb",  x"3c",  x"1f", -- 07D8
         x"fe",  x"28",  x"30",  x"11",  x"f6",  x"80",  x"67",  x"3e", -- 07E0
         x"ff",  x"82",  x"38",  x"09",  x"ab",  x"6f",  x"3a",  x"d6", -- 07E8
         x"b7",  x"57",  x"0a",  x"c1",  x"c9",  x"c1",  x"37",  x"c9", -- 07F0
         x"7f",  x"7f",  x"44",  x"20",  x"03",  x"fe",  x"03",  x"30", -- 07F8
         x"08",  x"0e",  x"08",  x"fe",  x"02",  x"30",  x"02",  x"1e", -- 0800
         x"04",  x"d5",  x"cd",  x"a6",  x"d7",  x"cd",  x"db",  x"f4", -- 0808
         x"cd",  x"7c",  x"e3",  x"38",  x"06",  x"1d",  x"20",  x"f2", -- 0810
         x"cd",  x"f0",  x"f3",  x"d1",  x"fe",  x"03",  x"c8",  x"fe", -- 0818
         x"0f",  x"20",  x"05",  x"cd",  x"d5",  x"f3",  x"18",  x"f0", -- 0820
         x"fe",  x"13",  x"20",  x"dd",  x"18",  x"07",  x"4b",  x"fe", -- 0828
         x"02",  x"30",  x"02",  x"0e",  x"01",  x"cd",  x"a6",  x"d7", -- 0830
         x"3e",  x"05",  x"32",  x"a0",  x"b7",  x"cd",  x"99",  x"f4", -- 0838
         x"d8",  x"e5",  x"cd",  x"eb",  x"f4",  x"7e",  x"e1",  x"38", -- 0840
         x"56",  x"a7",  x"28",  x"e9",  x"2a",  x"97",  x"b7",  x"e5", -- 0848
         x"cd",  x"eb",  x"f4",  x"7e",  x"a7",  x"23",  x"7e",  x"e1", -- 0850
         x"28",  x"04",  x"cd",  x"70",  x"fb",  x"23",  x"1a",  x"fe", -- 0858
         x"2e",  x"c8",  x"fe",  x"2c",  x"20",  x"05",  x"13",  x"1a", -- 0860
         x"13",  x"18",  x"ef",  x"fe",  x"3a",  x"20",  x"06",  x"06", -- 0868
         x"00",  x"ed",  x"42",  x"18",  x"c0",  x"fe",  x"2f",  x"20", -- 0870
         x"0b",  x"13",  x"cd",  x"eb",  x"f4",  x"38",  x"20",  x"2a", -- 0878
         x"97",  x"b7",  x"18",  x"b1",  x"fe",  x"27",  x"20",  x"10", -- 0880
         x"13",  x"1a",  x"13",  x"a7",  x"28",  x"a7",  x"fe",  x"27", -- 0888
         x"28",  x"cc",  x"cd",  x"70",  x"fb",  x"23",  x"18",  x"f1", -- 0890
         x"a7",  x"28",  x"9a",  x"fe",  x"20",  x"28",  x"b0",  x"cd", -- 0898
         x"d1",  x"f4",  x"18",  x"91",  x"cd",  x"ff",  x"f5",  x"cd", -- 08A0
         x"ef",  x"c8",  x"da",  x"d1",  x"f4",  x"3e",  x"0d",  x"cd", -- 08A8
         x"e9",  x"b7",  x"3e",  x"0a",  x"c3",  x"e9",  x"b7",  x"3a", -- 08B0
         x"e1",  x"b7",  x"e6",  x"f0",  x"0f",  x"0f",  x"0f",  x"18", -- 08B8
         x"3d",  x"cd",  x"5c",  x"c9",  x"af",  x"d3",  x"91",  x"db", -- 08C0
         x"91",  x"c6",  x"ff",  x"d8",  x"c5",  x"21",  x"11",  x"fa", -- 08C8
         x"18",  x"57",  x"2e",  x"07",  x"cd",  x"52",  x"c9",  x"c5", -- 08D0
         x"45",  x"cd",  x"8a",  x"c3",  x"50",  x"38",  x"70",  x"3a", -- 08D8
         x"e4",  x"b7",  x"47",  x"2a",  x"e2",  x"b7",  x"7b",  x"cd", -- 08E0
         x"da",  x"c9",  x"21",  x"29",  x"fa",  x"18",  x"3a",  x"67", -- 08E8
         x"3e",  x"05",  x"bc",  x"d8",  x"20",  x"c1",  x"3a",  x"8a", -- 08F0
         x"b7",  x"fe",  x"0d",  x"30",  x"53",  x"87",  x"57",  x"7c", -- 08F8
         x"a7",  x"28",  x"cf",  x"7d",  x"a7",  x"28",  x"ba",  x"c5", -- 0900
         x"45",  x"0e",  x"80",  x"ed",  x"78",  x"c1",  x"d6",  x"ee", -- 0908
         x"28",  x"c2",  x"3d",  x"20",  x"3b",  x"cd",  x"5c",  x"c9", -- 0910
         x"c5",  x"3e",  x"02",  x"16",  x"01",  x"cd",  x"9c",  x"c3", -- 0918
         x"21",  x"4d",  x"d9",  x"cd",  x"0d",  x"ca",  x"21",  x"00", -- 0920
         x"fa",  x"22",  x"ea",  x"b7",  x"e1",  x"22",  x"99",  x"b7", -- 0928
         x"7b",  x"32",  x"e1",  x"b7",  x"21",  x"ef",  x"f9",  x"01", -- 0930
         x"bf",  x"f4",  x"a7",  x"cb",  x"4b",  x"20",  x"08",  x"22", -- 0938
         x"be",  x"b7",  x"ed",  x"43",  x"c1",  x"b7",  x"c9",  x"22", -- 0940
         x"c4",  x"b7",  x"ed",  x"43",  x"c7",  x"b7",  x"c9",  x"e1", -- 0948
         x"37",  x"c9",  x"3e",  x"01",  x"bc",  x"30",  x"05",  x"1d", -- 0950
         x"93",  x"38",  x"f4",  x"bb",  x"5a",  x"cb",  x"13",  x"3e", -- 0958
         x"02",  x"57",  x"bc",  x"30",  x"06",  x"79",  x"92",  x"ba", -- 0960
         x"30",  x"e5",  x"0f",  x"cb",  x"13",  x"01",  x"bf",  x"f4", -- 0968
         x"14",  x"7a",  x"bc",  x"30",  x"0d",  x"3a",  x"88",  x"b7", -- 0970
         x"a7",  x"28",  x"07",  x"92",  x"30",  x"d1",  x"01",  x"c2", -- 0978
         x"f9",  x"0f",  x"cb",  x"13",  x"c9",  x"cd",  x"ff",  x"f5", -- 0980
         x"67",  x"3e",  x"03",  x"bc",  x"d8",  x"16",  x"00",  x"cd", -- 0988
         x"52",  x"c9",  x"e5",  x"3a",  x"e7",  x"b7",  x"47",  x"2a", -- 0990
         x"e5",  x"b7",  x"23",  x"18",  x"17",  x"3e",  x"80",  x"18", -- 0998
         x"10",  x"7e",  x"e6",  x"07",  x"28",  x"11",  x"23",  x"fe", -- 09A0
         x"03",  x"28",  x"f2",  x"fe",  x"05",  x"20",  x"05",  x"3e", -- 09A8
         x"68",  x"a6",  x"b3",  x"5f",  x"05",  x"28",  x"98",  x"23", -- 09B0
         x"10",  x"e7",  x"e1",  x"7c",  x"06",  x"07",  x"a7",  x"28", -- 09B8
         x"01",  x"45",  x"cd",  x"8a",  x"c3",  x"d8",  x"21",  x"41", -- 09C0
         x"fa",  x"01",  x"4c",  x"fa",  x"cd",  x"3b",  x"c9",  x"3a", -- 09C8
         x"e7",  x"b7",  x"47",  x"2a",  x"e5",  x"b7",  x"7b",  x"32", -- 09D0
         x"e8",  x"b7",  x"e6",  x"04",  x"0f",  x"0f",  x"c6",  x"0c", -- 09D8
         x"4f",  x"78",  x"06",  x"02",  x"90",  x"f3",  x"ed",  x"b3", -- 09E0
         x"47",  x"0d",  x"0d",  x"ed",  x"b3",  x"fb",  x"a7",  x"c9", -- 09E8
         x"21",  x"24",  x"d8",  x"11",  x"00",  x"a8",  x"01",  x"12", -- 09F0
         x"00",  x"ed",  x"b0",  x"af",  x"cd",  x"ef",  x"c8",  x"d8", -- 09F8
         x"7a",  x"32",  x"00",  x"a8",  x"21",  x"41",  x"fa",  x"22", -- 0A00
         x"c4",  x"b7",  x"21",  x"36",  x"d8",  x"56",  x"23",  x"c3", -- 0A08
         x"61",  x"f5",  x"f5",  x"3a",  x"e1",  x"b7",  x"cb",  x"7f", -- 0A10
         x"28",  x"29",  x"e6",  x"f0",  x"fe",  x"90",  x"28",  x"17", -- 0A18
         x"fe",  x"a0",  x"20",  x"1f",  x"f1",  x"e5",  x"c5",  x"21", -- 0A20
         x"75",  x"d9",  x"01",  x"07",  x"00",  x"ed",  x"b1",  x"20", -- 0A28
         x"0f",  x"0e",  x"06",  x"09",  x"7e",  x"18",  x"09",  x"f1", -- 0A30
         x"fe",  x"7e",  x"20",  x"08",  x"3e",  x"83",  x"18",  x"04", -- 0A38
         x"c1",  x"e1",  x"f5",  x"f1",  x"fe",  x"09",  x"28",  x"0d", -- 0A40
         x"f5",  x"3a",  x"a2",  x"b7",  x"cb",  x"5f",  x"28",  x"0e", -- 0A48
         x"f1",  x"fe",  x"7f",  x"20",  x"02",  x"3e",  x"20",  x"fe", -- 0A50
         x"20",  x"30",  x"04",  x"3e",  x"5f",  x"f5",  x"f1",  x"c3", -- 0A58
         x"e9",  x"b7",  x"e5",  x"d5",  x"3a",  x"e1",  x"b7",  x"cb", -- 0A60
         x"47",  x"20",  x"2e",  x"2a",  x"b9",  x"b7",  x"5f",  x"7e", -- 0A68
         x"a7",  x"20",  x"12",  x"cb",  x"4b",  x"21",  x"ec",  x"f9", -- 0A70
         x"11",  x"0b",  x"f0",  x"20",  x"12",  x"11",  x"08",  x"f0", -- 0A78
         x"22",  x"be",  x"b7",  x"18",  x"0d",  x"21",  x"ef",  x"f9", -- 0A80
         x"11",  x"05",  x"f0",  x"fe",  x"02",  x"28",  x"f1",  x"22", -- 0A88
         x"c4",  x"b7",  x"ed",  x"53",  x"b9",  x"b7",  x"d1",  x"e1", -- 0A90
         x"c9",  x"c5",  x"f5",  x"e6",  x"f0",  x"f2",  x"c4",  x"ca", -- 0A98
         x"2a",  x"cb",  x"b7",  x"06",  x"20",  x"0e",  x"28",  x"7e", -- 0AA0
         x"23",  x"fe",  x"20",  x"30",  x"02",  x"3e",  x"20",  x"cd", -- 0AA8
         x"ef",  x"f9",  x"0d",  x"20",  x"f2",  x"3e",  x"0d",  x"cd", -- 0AB0
         x"44",  x"ca",  x"3e",  x"0a",  x"cd",  x"44",  x"ca",  x"10", -- 0AB8
         x"e4",  x"c3",  x"97",  x"e0",  x"e6",  x"f0",  x"fe",  x"10", -- 0AC0
         x"ca",  x"92",  x"cb",  x"fe",  x"20",  x"ca",  x"d0",  x"cb", -- 0AC8
         x"fe",  x"30",  x"ca",  x"fe",  x"cb",  x"fe",  x"50",  x"28", -- 0AD0
         x"3b",  x"fe",  x"70",  x"28",  x"67",  x"26",  x"00",  x"cd", -- 0AD8
         x"9d",  x"cc",  x"2e",  x"00",  x"0e",  x"08",  x"cd",  x"c3", -- 0AE0
         x"cc",  x"e5",  x"06",  x"08",  x"21",  x"00",  x"b7",  x"cb", -- 0AE8
         x"16",  x"17",  x"23",  x"10",  x"fa",  x"cd",  x"e9",  x"b7", -- 0AF0
         x"0d",  x"20",  x"ef",  x"e1",  x"2c",  x"3e",  x"28",  x"bd", -- 0AF8
         x"20",  x"e2",  x"7c",  x"c6",  x"08",  x"67",  x"30",  x"d7", -- 0B00
         x"3e",  x"0d",  x"cd",  x"e9",  x"b7",  x"3e",  x"0a",  x"cd", -- 0B08
         x"e9",  x"b7",  x"18",  x"ad",  x"21",  x"00",  x"00",  x"cd", -- 0B10
         x"9d",  x"cc",  x"0e",  x"18",  x"cd",  x"c3",  x"cc",  x"cd", -- 0B18
         x"7e",  x"cc",  x"20",  x"f6",  x"7c",  x"c6",  x"18",  x"67", -- 0B20
         x"2e",  x"00",  x"fe",  x"f0",  x"20",  x"e9",  x"cd",  x"9d", -- 0B28
         x"cc",  x"0e",  x"10",  x"cd",  x"c3",  x"cc",  x"06",  x"08", -- 0B30
         x"af",  x"12",  x"13",  x"10",  x"fc",  x"cd",  x"7e",  x"cc", -- 0B38
         x"20",  x"ef",  x"18",  x"c4",  x"26",  x"00",  x"cd",  x"9d", -- 0B40
         x"cc",  x"2e",  x"00",  x"06",  x"08",  x"e5",  x"cd",  x"4c", -- 0B48
         x"e0",  x"11",  x"00",  x"b7",  x"7e",  x"12",  x"13",  x"12", -- 0B50
         x"13",  x"12",  x"13",  x"2c",  x"10",  x"f6",  x"0e",  x"08", -- 0B58
         x"06",  x"18",  x"21",  x"00",  x"b7",  x"cb",  x"16",  x"cb", -- 0B60
         x"13",  x"cb",  x"12",  x"17",  x"23",  x"10",  x"f6",  x"77", -- 0B68
         x"06",  x"03",  x"7e",  x"cd",  x"e9",  x"b7",  x"7a",  x"cd", -- 0B70
         x"e9",  x"b7",  x"7b",  x"cd",  x"e9",  x"b7",  x"10",  x"f2", -- 0B78
         x"0d",  x"20",  x"dd",  x"e1",  x"2c",  x"3e",  x"28",  x"bd", -- 0B80
         x"20",  x"c1",  x"7c",  x"c6",  x"08",  x"67",  x"30",  x"b6", -- 0B88
         x"18",  x"3b",  x"26",  x"00",  x"cd",  x"9d",  x"cc",  x"2e", -- 0B90
         x"00",  x"06",  x"04",  x"e5",  x"cd",  x"4c",  x"e0",  x"11", -- 0B98
         x"00",  x"b7",  x"7e",  x"12",  x"13",  x"12",  x"13",  x"2c", -- 0BA0
         x"10",  x"f8",  x"0e",  x"08",  x"06",  x"08",  x"21",  x"00", -- 0BA8
         x"b7",  x"cb",  x"16",  x"17",  x"23",  x"10",  x"fa",  x"cd", -- 0BB0
         x"e9",  x"b7",  x"cd",  x"e9",  x"b7",  x"0d",  x"20",  x"ec", -- 0BB8
         x"e1",  x"2c",  x"3e",  x"28",  x"bd",  x"20",  x"d2",  x"7c", -- 0BC0
         x"c6",  x"04",  x"67",  x"30",  x"c7",  x"c3",  x"08",  x"cb", -- 0BC8
         x"cd",  x"9d",  x"cc",  x"06",  x"2a",  x"21",  x"00",  x"00", -- 0BD0
         x"0e",  x"06",  x"cd",  x"c3",  x"cc",  x"cd",  x"2a",  x"cc", -- 0BD8
         x"20",  x"f6",  x"3e",  x"06",  x"84",  x"67",  x"2e",  x"00", -- 0BE0
         x"cd",  x"9d",  x"cc",  x"05",  x"20",  x"ea",  x"0e",  x"04", -- 0BE8
         x"cd",  x"c3",  x"cc",  x"af",  x"12",  x"13",  x"12",  x"cd", -- 0BF0
         x"2a",  x"cc",  x"20",  x"f2",  x"18",  x"cf",  x"cd",  x"9d", -- 0BF8
         x"cc",  x"06",  x"55",  x"21",  x"00",  x"00",  x"0e",  x"03", -- 0C00
         x"cd",  x"d1",  x"cc",  x"cd",  x"53",  x"cc",  x"20",  x"f6", -- 0C08
         x"24",  x"24",  x"24",  x"2e",  x"00",  x"cd",  x"9d",  x"cc", -- 0C10
         x"10",  x"ec",  x"0e",  x"04",  x"cd",  x"d1",  x"cc",  x"af", -- 0C18
         x"12",  x"13",  x"12",  x"cd",  x"53",  x"cc",  x"20",  x"f2", -- 0C20
         x"18",  x"a3",  x"e5",  x"c5",  x"2e",  x"80",  x"06",  x"00", -- 0C28
         x"11",  x"00",  x"b7",  x"1a",  x"a5",  x"28",  x"01",  x"37", -- 0C30
         x"cb",  x"10",  x"13",  x"3e",  x"06",  x"bb",  x"20",  x"f3", -- 0C38
         x"a7",  x"cb",  x"10",  x"78",  x"cd",  x"e9",  x"b7",  x"cb", -- 0C40
         x"0d",  x"f2",  x"2e",  x"cc",  x"c1",  x"e1",  x"2c",  x"3e", -- 0C48
         x"28",  x"bd",  x"c9",  x"e5",  x"c5",  x"2e",  x"80",  x"06", -- 0C50
         x"00",  x"11",  x"00",  x"b7",  x"1a",  x"a5",  x"28",  x"01", -- 0C58
         x"37",  x"cb",  x"10",  x"13",  x"3e",  x"06",  x"bb",  x"20", -- 0C60
         x"f3",  x"78",  x"17",  x"17",  x"cd",  x"e9",  x"b7",  x"cd", -- 0C68
         x"e9",  x"b7",  x"cb",  x"0d",  x"f2",  x"57",  x"cc",  x"c1", -- 0C70
         x"e1",  x"2c",  x"3e",  x"28",  x"bd",  x"c9",  x"e5",  x"1e", -- 0C78
         x"08",  x"0e",  x"03",  x"21",  x"00",  x"b7",  x"06",  x"08", -- 0C80
         x"cb",  x"16",  x"17",  x"23",  x"10",  x"fa",  x"cd",  x"e9", -- 0C88
         x"b7",  x"0d",  x"20",  x"f2",  x"1d",  x"20",  x"ea",  x"e1", -- 0C90
         x"2c",  x"3e",  x"28",  x"bd",  x"c9",  x"e5",  x"c5",  x"af", -- 0C98
         x"21",  x"e1",  x"b7",  x"ed",  x"6f",  x"4f",  x"ed",  x"67", -- 0CA0
         x"0c",  x"21",  x"c5",  x"d7",  x"46",  x"0d",  x"28",  x"09", -- 0CA8
         x"04",  x"7d",  x"80",  x"6f",  x"30",  x"f6",  x"24",  x"18", -- 0CB0
         x"f3",  x"23",  x"7e",  x"cd",  x"e9",  x"b7",  x"10",  x"f9", -- 0CB8
         x"c1",  x"e1",  x"c9",  x"e5",  x"c5",  x"cd",  x"4c",  x"e0", -- 0CC0
         x"11",  x"00",  x"b7",  x"06",  x"00",  x"ed",  x"b0",  x"18", -- 0CC8
         x"ef",  x"e5",  x"cd",  x"4c",  x"e0",  x"11",  x"00",  x"b7", -- 0CD0
         x"7e",  x"12",  x"13",  x"12",  x"13",  x"2c",  x"0d",  x"20", -- 0CD8
         x"f7",  x"e1",  x"c9",  x"5a",  x"57",  x"d5",  x"c5",  x"cb", -- 0CE0
         x"5b",  x"28",  x"32",  x"dd",  x"cb",  x"07",  x"ce",  x"3e", -- 0CE8
         x"d5",  x"be",  x"d5",  x"11",  x"a0",  x"00",  x"20",  x"03", -- 0CF0
         x"11",  x"00",  x"05",  x"ed",  x"53",  x"d8",  x"b7",  x"cd", -- 0CF8
         x"8a",  x"d7",  x"11",  x"00",  x"b7",  x"cd",  x"97",  x"ed", -- 0D00
         x"20",  x"05",  x"01",  x"0b",  x"00",  x"ed",  x"b0",  x"eb", -- 0D08
         x"d1",  x"72",  x"2c",  x"7d",  x"32",  x"da",  x"b7",  x"a7", -- 0D10
         x"c1",  x"d1",  x"cb",  x"9b",  x"c9",  x"2a",  x"da",  x"b7", -- 0D18
         x"26",  x"b7",  x"72",  x"cb",  x"73",  x"20",  x"26",  x"2c", -- 0D20
         x"f2",  x"13",  x"cd",  x"dd",  x"cb",  x"07",  x"4e",  x"20", -- 0D28
         x"08",  x"cd",  x"5e",  x"ce",  x"38",  x"e2",  x"af",  x"18", -- 0D30
         x"db",  x"dd",  x"cb",  x"07",  x"8e",  x"21",  x"f5",  x"b7", -- 0D38
         x"cd",  x"c9",  x"e4",  x"02",  x"38",  x"d2",  x"cd",  x"6a", -- 0D40
         x"ce",  x"38",  x"cd",  x"18",  x"e9",  x"dd",  x"cb",  x"07", -- 0D48
         x"4e",  x"28",  x"09",  x"21",  x"f5",  x"b7",  x"cd",  x"c9", -- 0D50
         x"e4",  x"02",  x"18",  x"04",  x"cd",  x"5e",  x"ce",  x"d8", -- 0D58
         x"ed",  x"4b",  x"d8",  x"b7",  x"cd",  x"c9",  x"e4",  x"03", -- 0D60
         x"f5",  x"cd",  x"db",  x"f4",  x"f1",  x"18",  x"a9",  x"cd", -- 0D68
         x"c9",  x"e4",  x"05",  x"dd",  x"cb",  x"07",  x"ae",  x"18", -- 0D70
         x"9f",  x"5a",  x"d5",  x"c5",  x"cb",  x"73",  x"20",  x"ef", -- 0D78
         x"cb",  x"5b",  x"28",  x"67",  x"e5",  x"cd",  x"8a",  x"d7", -- 0D80
         x"21",  x"f5",  x"b7",  x"cd",  x"c9",  x"e4",  x"04",  x"e1", -- 0D88
         x"da",  x"46",  x"ce",  x"dd",  x"7e",  x"02",  x"fe",  x"01", -- 0D90
         x"c2",  x"46",  x"ce",  x"dd",  x"cb",  x"07",  x"be",  x"dd", -- 0D98
         x"34",  x"03",  x"11",  x"00",  x"b7",  x"cd",  x"97",  x"ed", -- 0DA0
         x"20",  x"36",  x"06",  x"0b",  x"1a",  x"fe",  x"d5",  x"20", -- 0DA8
         x"04",  x"dd",  x"cb",  x"07",  x"ee",  x"c6",  x"29",  x"30", -- 0DB0
         x"0d",  x"1a",  x"d6",  x"04",  x"12",  x"13",  x"12",  x"13", -- 0DB8
         x"12",  x"32",  x"5e",  x"03",  x"1b",  x"1b",  x"1a",  x"cd", -- 0DC0
         x"8c",  x"e0",  x"be",  x"28",  x"04",  x"dd",  x"cb",  x"07", -- 0DC8
         x"fe",  x"23",  x"13",  x"10",  x"f1",  x"cd",  x"db",  x"f4", -- 0DD0
         x"dd",  x"cb",  x"07",  x"7e",  x"37",  x"c2",  x"18",  x"cd", -- 0DD8
         x"eb",  x"56",  x"2c",  x"7d",  x"32",  x"da",  x"b7",  x"7a", -- 0DE0
         x"c3",  x"17",  x"cd",  x"2a",  x"da",  x"b7",  x"26",  x"b7", -- 0DE8
         x"cb",  x"7d",  x"28",  x"ed",  x"cd",  x"c9",  x"e4",  x"01", -- 0DF0
         x"38",  x"36",  x"3e",  x"ff",  x"dd",  x"be",  x"02",  x"28", -- 0DF8
         x"1a",  x"dd",  x"7e",  x"03",  x"dd",  x"be",  x"02",  x"28", -- 0E00
         x"12",  x"3e",  x"2a",  x"cd",  x"8c",  x"e0",  x"cd",  x"c9", -- 0E08
         x"f0",  x"19",  x"00",  x"cd",  x"7c",  x"e3",  x"30",  x"dc", -- 0E10
         x"c3",  x"18",  x"cd",  x"dd",  x"34",  x"03",  x"3d",  x"dd", -- 0E18
         x"cb",  x"07",  x"6e",  x"20",  x"06",  x"cd",  x"c9",  x"f0", -- 0E20
         x"3e",  x"19",  x"00",  x"21",  x"00",  x"b7",  x"18",  x"b1", -- 0E28
         x"cd",  x"97",  x"ed",  x"20",  x"14",  x"cd",  x"cf",  x"f0", -- 0E30
         x"09",  x"09",  x"09",  x"09",  x"3f",  x"00",  x"cd",  x"c9", -- 0E38
         x"f0",  x"0d",  x"0a",  x"00",  x"18",  x"cd",  x"cd",  x"97", -- 0E40
         x"ed",  x"37",  x"20",  x"cc",  x"cd",  x"cf",  x"f0",  x"2a", -- 0E48
         x"08",  x"00",  x"cd",  x"7c",  x"e3",  x"38",  x"c1",  x"cd", -- 0E50
         x"c9",  x"e4",  x"01",  x"c3",  x"90",  x"cd",  x"ed",  x"4b", -- 0E58
         x"d8",  x"b7",  x"cd",  x"c9",  x"e4",  x"00",  x"d8",  x"cd", -- 0E60
         x"c0",  x"e4",  x"cd",  x"c9",  x"f0",  x"19",  x"00",  x"c3", -- 0E68
         x"7c",  x"e3",  x"00",  x"56",  x"41",  x"52",  x"49",  x"41", -- 0E70
         x"42",  x"45",  x"4c",  x"00",  x"01",  x"53",  x"54",  x"41", -- 0E78
         x"52",  x"54",  x"2d",  x"52",  x"4f",  x"4d",  x"00",  x"70", -- 0E80
         x"33",  x"32",  x"4b",  x"20",  x"45",  x"50",  x"52",  x"4f", -- 0E88
         x"4d",  x"00",  x"71",  x"36",  x"34",  x"4b",  x"20",  x"45", -- 0E90
         x"50",  x"52",  x"4f",  x"4d",  x"00",  x"72",  x"31",  x"32", -- 0E98
         x"38",  x"4b",  x"20",  x"45",  x"50",  x"52",  x"4f",  x"4d", -- 0EA0
         x"00",  x"73",  x"32",  x"35",  x"36",  x"4b",  x"20",  x"45", -- 0EA8
         x"50",  x"52",  x"4f",  x"4d",  x"00",  x"77",  x"36",  x"34", -- 0EB0
         x"4b",  x"20",  x"52",  x"41",  x"4d",  x"00",  x"78",  x"31", -- 0EB8
         x"32",  x"38",  x"4b",  x"20",  x"52",  x"41",  x"4d",  x"00", -- 0EC0
         x"79",  x"32",  x"35",  x"36",  x"4b",  x"20",  x"52",  x"41", -- 0EC8
         x"4d",  x"00",  x"7a",  x"35",  x"31",  x"32",  x"4b",  x"20", -- 0ED0
         x"52",  x"41",  x"4d",  x"00",  x"7b",  x"31",  x"4d",  x"20", -- 0ED8
         x"52",  x"41",  x"4d",  x"00",  x"a7",  x"46",  x"4c",  x"4f", -- 0EE0
         x"50",  x"50",  x"59",  x"00",  x"d9",  x"45",  x"50",  x"52", -- 0EE8
         x"4f",  x"4d",  x"4d",  x"45",  x"52",  x"20",  x"33",  x"32", -- 0EF0
         x"4b",  x"00",  x"da",  x"50",  x"49",  x"4f",  x"2d",  x"33", -- 0EF8
         x"00",  x"db",  x"45",  x"50",  x"52",  x"4f",  x"4d",  x"4d", -- 0F00
         x"45",  x"52",  x"20",  x"36",  x"34",  x"4b",  x"00",  x"dc", -- 0F08
         x"53",  x"4f",  x"55",  x"4e",  x"44",  x"00",  x"e3",  x"44", -- 0F10
         x"41",  x"55",  x"31",  x"00",  x"e7",  x"41",  x"44",  x"55", -- 0F18
         x"31",  x"00",  x"ec",  x"53",  x"43",  x"41",  x"4e",  x"4e", -- 0F20
         x"45",  x"52",  x"00",  x"ee",  x"56",  x"2e",  x"32",  x"34", -- 0F28
         x"00",  x"ef",  x"44",  x"49",  x"47",  x"49",  x"54",  x"41", -- 0F30
         x"4c",  x"20",  x"49",  x"2f",  x"4f",  x"00",  x"f0",  x"38", -- 0F38
         x"4b",  x"20",  x"43",  x"4d",  x"4f",  x"53",  x"2d",  x"52", -- 0F40
         x"41",  x"4d",  x"00",  x"f1",  x"31",  x"36",  x"4b",  x"20", -- 0F48
         x"43",  x"4d",  x"4f",  x"53",  x"2d",  x"52",  x"41",  x"4d", -- 0F50
         x"00",  x"f2",  x"33",  x"32",  x"4b",  x"20",  x"43",  x"4d", -- 0F58
         x"4f",  x"53",  x"2d",  x"52",  x"41",  x"4d",  x"00",  x"f4", -- 0F60
         x"31",  x"36",  x"4b",  x"20",  x"52",  x"41",  x"4d",  x"00", -- 0F68
         x"f5",  x"33",  x"32",  x"4b",  x"20",  x"52",  x"41",  x"4d", -- 0F70
         x"00",  x"f6",  x"36",  x"34",  x"4b",  x"20",  x"52",  x"41", -- 0F78
         x"4d",  x"00",  x"f7",  x"38",  x"4b",  x"20",  x"52",  x"4f", -- 0F80
         x"4d",  x"00",  x"f8",  x"31",  x"36",  x"4b",  x"20",  x"52", -- 0F88
         x"4f",  x"4d",  x"00",  x"f9",  x"47",  x"49",  x"44",  x"45", -- 0F90
         x"00",  x"fc",  x"42",  x"41",  x"53",  x"49",  x"43",  x"00", -- 0F98
         x"ff",  x"3f",  x"3f",  x"3f",  x"00",  x"53",  x"4f",  x"46", -- 0FA0
         x"54",  x"57",  x"41",  x"52",  x"45",  x"00",  x"55",  x"53", -- 0FA8
         x"45",  x"52",  x"00",  x"4e",  x"45",  x"54",  x"2b",  x"55", -- 0FB0
         x"53",  x"42",  x"00",  x"34",  x"2a",  x"38",  x"4b",  x"20", -- 0FB8
         x"52",  x"41",  x"4d",  x"00",  x"38",  x"2a",  x"38",  x"4b", -- 0FC0
         x"20",  x"45",  x"50",  x"52",  x"4f",  x"4d",  x"00",  x"ff", -- 0FC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FF8
         x"f3",  x"db",  x"88",  x"f6",  x"60",  x"cd",  x"58",  x"e4", -- 1000
         x"dd",  x"36",  x"02",  x"00",  x"01",  x"00",  x"10",  x"dd", -- 1008
         x"34",  x"02",  x"3e",  x"87",  x"f3",  x"d3",  x"8d",  x"3e", -- 1010
         x"2f",  x"d3",  x"8d",  x"fb",  x"5f",  x"cd",  x"62",  x"d0", -- 1018
         x"ed",  x"a1",  x"ea",  x"1d",  x"d0",  x"cd",  x"60",  x"d0", -- 1020
         x"dd",  x"7e",  x"02",  x"cd",  x"4d",  x"d0",  x"dd",  x"6e", -- 1028
         x"05",  x"dd",  x"66",  x"06",  x"06",  x"80",  x"7e",  x"cd", -- 1030
         x"4d",  x"d0",  x"79",  x"86",  x"4f",  x"23",  x"10",  x"f6", -- 1038
         x"cd",  x"4d",  x"d0",  x"cd",  x"65",  x"d0",  x"5d",  x"54", -- 1040
         x"3e",  x"03",  x"d3",  x"8d",  x"c9",  x"c5",  x"4f",  x"06", -- 1048
         x"08",  x"cb",  x"09",  x"1e",  x"17",  x"d4",  x"62",  x"d0", -- 1050
         x"1e",  x"2f",  x"dc",  x"62",  x"d0",  x"10",  x"f2",  x"c1", -- 1058
         x"1e",  x"5d",  x"cd",  x"65",  x"d0",  x"dd",  x"73",  x"00", -- 1060
         x"dd",  x"7e",  x"00",  x"a7",  x"20",  x"fa",  x"c9",  x"cd", -- 1068
         x"4d",  x"e4",  x"3e",  x"83",  x"d3",  x"8a",  x"e5",  x"d5", -- 1070
         x"06",  x"16",  x"cd",  x"cd",  x"d0",  x"38",  x"f9",  x"fe", -- 1078
         x"ba",  x"cd",  x"c2",  x"d0",  x"38",  x"f2",  x"10",  x"f2", -- 1080
         x"06",  x"02",  x"af",  x"cd",  x"d1",  x"d0",  x"fe",  x"5d", -- 1088
         x"30",  x"f6",  x"10",  x"f6",  x"dd",  x"6e",  x"05",  x"dd", -- 1090
         x"66",  x"06",  x"cd",  x"e2",  x"d0",  x"38",  x"1b",  x"dd", -- 1098
         x"77",  x"02",  x"06",  x"80",  x"1e",  x"00",  x"cd",  x"e2", -- 10A0
         x"d0",  x"38",  x"0f",  x"77",  x"83",  x"5f",  x"23",  x"10", -- 10A8
         x"f5",  x"6f",  x"cd",  x"e2",  x"d0",  x"38",  x"03",  x"95", -- 10B0
         x"c6",  x"ff",  x"d1",  x"e1",  x"f3",  x"3e",  x"03",  x"d3", -- 10B8
         x"8a",  x"fb",  x"db",  x"88",  x"cb",  x"ef",  x"30",  x"02", -- 10C0
         x"cb",  x"af",  x"d3",  x"88",  x"c9",  x"af",  x"cd",  x"d1", -- 10C8
         x"d0",  x"4f",  x"dd",  x"36",  x"00",  x"00",  x"db",  x"88", -- 10D0
         x"d3",  x"88",  x"af",  x"dd",  x"b6",  x"00",  x"28",  x"f6", -- 10D8
         x"81",  x"c9",  x"16",  x"80",  x"cd",  x"cd",  x"d0",  x"38", -- 10E0
         x"03",  x"fe",  x"ba",  x"d8",  x"3f",  x"cb",  x"1a",  x"30", -- 10E8
         x"f3",  x"cd",  x"cd",  x"d0",  x"7a",  x"c9",  x"dd",  x"36", -- 10F0
         x"02",  x"00",  x"dd",  x"36",  x"03",  x"01",  x"cd",  x"94", -- 10F8
         x"d1",  x"3e",  x"09",  x"21",  x"3e",  x"01",  x"cd",  x"4a", -- 1100
         x"d1",  x"d8",  x"0d",  x"e5",  x"dd",  x"6e",  x"05",  x"dd", -- 1108
         x"66",  x"06",  x"ed",  x"78",  x"cd",  x"70",  x"fb",  x"23", -- 1110
         x"04",  x"20",  x"f7",  x"e1",  x"dd",  x"34",  x"02",  x"c9", -- 1118
         x"3e",  x"41",  x"18",  x"26",  x"dd",  x"36",  x"02",  x"00", -- 1120
         x"cd",  x"94",  x"d1",  x"3e",  x"0b",  x"21",  x"3e",  x"03", -- 1128
         x"dd",  x"34",  x"02",  x"dd",  x"6e",  x"05",  x"dd",  x"66", -- 1130
         x"06",  x"01",  x"f2",  x"80",  x"1e",  x"80",  x"08",  x"cd", -- 1138
         x"80",  x"fb",  x"ed",  x"79",  x"23",  x"04",  x"1d",  x"20", -- 1140
         x"f6",  x"08",  x"01",  x"f3",  x"80",  x"ed",  x"79",  x"c5", -- 1148
         x"3e",  x"01",  x"cd",  x"a3",  x"e2",  x"c1",  x"ed",  x"78", -- 1150
         x"a7",  x"cb",  x"47",  x"20",  x"f2",  x"cb",  x"7f",  x"c8", -- 1158
         x"01",  x"f1",  x"83",  x"ed",  x"78",  x"fe",  x"20",  x"30", -- 1160
         x"0d",  x"01",  x"f3",  x"81",  x"ed",  x"78",  x"cd",  x"c4", -- 1168
         x"f3",  x"cd",  x"d1",  x"f4",  x"37",  x"c9",  x"06",  x"00", -- 1170
         x"ed",  x"78",  x"04",  x"a7",  x"28",  x"f6",  x"cd",  x"d5", -- 1178
         x"f3",  x"18",  x"f5",  x"01",  x"f1",  x"80",  x"18",  x"c5", -- 1180
         x"dd",  x"36",  x"02",  x"fe",  x"cd",  x"2e",  x"d1",  x"d8", -- 1188
         x"3e",  x"43",  x"18",  x"b6",  x"11",  x"0c",  x"ff",  x"01", -- 1190
         x"f3",  x"82",  x"7e",  x"ed",  x"79",  x"a2",  x"28",  x"01", -- 1198
         x"23",  x"04",  x"1d",  x"20",  x"f5",  x"c9",  x"cd",  x"6a", -- 11A0
         x"f5",  x"d8",  x"11",  x"0c",  x"df",  x"cd",  x"97",  x"d1", -- 11A8
         x"eb",  x"13",  x"c9",  x"79",  x"01",  x"00",  x"dc",  x"87", -- 11B0
         x"38",  x"2c",  x"05",  x"fe",  x"40",  x"38",  x"27",  x"06", -- 11B8
         x"ed",  x"fe",  x"b6",  x"38",  x"21",  x"fe",  x"bc",  x"38", -- 11C0
         x"0c",  x"fe",  x"c0",  x"38",  x"19",  x"28",  x"06",  x"06", -- 11C8
         x"fc",  x"fe",  x"f6",  x"38",  x"11",  x"01",  x"b8",  x"da", -- 11D0
         x"d6",  x"b6",  x"fe",  x"06",  x"38",  x"08",  x"d6",  x"04", -- 11D8
         x"fe",  x"06",  x"28",  x"02",  x"d6",  x"34",  x"6f",  x"26", -- 11E0
         x"00",  x"29",  x"c3",  x"cb",  x"e0",  x"e5",  x"d5",  x"c5", -- 11E8
         x"f5",  x"08",  x"f5",  x"79",  x"08",  x"3a",  x"9e",  x"b7", -- 11F0
         x"e5",  x"d5",  x"ed",  x"a0",  x"ed",  x"a0",  x"ed",  x"a0", -- 11F8
         x"ed",  x"a0",  x"ed",  x"a0",  x"ed",  x"a0",  x"ed",  x"a0", -- 1200
         x"ed",  x"a0",  x"ea",  x"fa",  x"d1",  x"d1",  x"e1",  x"24", -- 1208
         x"14",  x"08",  x"4f",  x"08",  x"3d",  x"20",  x"e1",  x"08", -- 1210
         x"f1",  x"08",  x"c3",  x"97",  x"e0",  x"41",  x"55",  x"77", -- 1218
         x"2c",  x"77",  x"2c",  x"77",  x"2c",  x"77",  x"2c",  x"77", -- 1220
         x"2c",  x"77",  x"2c",  x"77",  x"2c",  x"77",  x"6a",  x"24", -- 1228
         x"10",  x"ec",  x"c9",  x"3a",  x"9e",  x"b7",  x"4f",  x"06", -- 1230
         x"00",  x"3a",  x"9f",  x"b7",  x"3d",  x"28",  x"3a",  x"d5", -- 1238
         x"f5",  x"50",  x"58",  x"cd",  x"68",  x"e0",  x"eb",  x"21", -- 1240
         x"28",  x"00",  x"19",  x"e5",  x"c5",  x"ed",  x"b0",  x"c1", -- 1248
         x"d1",  x"3d",  x"20",  x"f3",  x"f1",  x"87",  x"87",  x"87", -- 1250
         x"4f",  x"50",  x"58",  x"cd",  x"42",  x"e0",  x"eb",  x"2e", -- 1258
         x"08",  x"19",  x"3a",  x"a2",  x"b7",  x"1f",  x"1f",  x"38", -- 1260
         x"0b",  x"f5",  x"cd",  x"87",  x"f9",  x"cd",  x"ed",  x"d1", -- 1268
         x"cd",  x"87",  x"f9",  x"f1",  x"17",  x"d4",  x"ed",  x"d1", -- 1270
         x"d1",  x"15",  x"1e",  x"00",  x"cd",  x"68",  x"e0",  x"d8", -- 1278
         x"3a",  x"9e",  x"b7",  x"47",  x"4f",  x"af",  x"77",  x"23", -- 1280
         x"10",  x"fc",  x"cd",  x"42",  x"e0",  x"d8",  x"d5",  x"dd", -- 1288
         x"cb",  x"01",  x"5e",  x"3a",  x"a2",  x"b7",  x"20",  x"04", -- 1290
         x"cb",  x"77",  x"20",  x"1c",  x"0f",  x"5f",  x"38",  x"06", -- 1298
         x"af",  x"e5",  x"cd",  x"1d",  x"d2",  x"e1",  x"cb",  x"0b", -- 12A0
         x"38",  x"0c",  x"cd",  x"87",  x"f9",  x"3a",  x"a3",  x"b7", -- 12A8
         x"cd",  x"1d",  x"d2",  x"cd",  x"87",  x"f9",  x"d1",  x"c9", -- 12B0
         x"3a",  x"a3",  x"b7",  x"e6",  x"03",  x"1f",  x"3d",  x"2f", -- 12B8
         x"5f",  x"9f",  x"e5",  x"cd",  x"1d",  x"d2",  x"e1",  x"cd", -- 12C0
         x"87",  x"f9",  x"7b",  x"18",  x"e3",  x"af",  x"3d",  x"5f", -- 12C8
         x"57",  x"3c",  x"13",  x"13",  x"ed",  x"52",  x"30",  x"f9", -- 12D0
         x"c3",  x"9c",  x"fb",  x"af",  x"06",  x"08",  x"cb",  x"1a", -- 12D8
         x"30",  x"01",  x"81",  x"1f",  x"cb",  x"1a",  x"10",  x"f8", -- 12E0
         x"47",  x"7a",  x"c9",  x"7f",  x"7f",  x"76",  x"69",  x"65", -- 12E8
         x"77",  x"03",  x"7d",  x"fe",  x"10",  x"30",  x"0c",  x"7c", -- 12F0
         x"a7",  x"20",  x"08",  x"21",  x"82",  x"b7",  x"ed",  x"6f", -- 12F8
         x"66",  x"2e",  x"00",  x"11",  x"00",  x"88",  x"01",  x"00", -- 1300
         x"20",  x"cd",  x"80",  x"fb",  x"12",  x"23",  x"13",  x"0d", -- 1308
         x"20",  x"f7",  x"10",  x"f5",  x"3e",  x"0b",  x"cd",  x"8c", -- 1310
         x"e0",  x"3e",  x"08",  x"32",  x"a0",  x"b7",  x"cd",  x"21", -- 1318
         x"d3",  x"3e",  x"01",  x"4f",  x"cd",  x"c4",  x"f3",  x"79", -- 1320
         x"c6",  x"22",  x"30",  x"f7",  x"c9",  x"28",  x"14",  x"f5", -- 1328
         x"cd",  x"cf",  x"f0",  x"20",  x"4f",  x"4e",  x"00",  x"f1", -- 1330
         x"3e",  x"20",  x"30",  x"02",  x"3e",  x"2a",  x"cd",  x"d5", -- 1338
         x"f3",  x"18",  x"08",  x"cd",  x"cf",  x"f0",  x"20",  x"4f", -- 1340
         x"46",  x"46",  x"00",  x"c3",  x"db",  x"f4",  x"7d",  x"cd", -- 1348
         x"b9",  x"f3",  x"7c",  x"cd",  x"b9",  x"f3",  x"7a",  x"c3", -- 1350
         x"b9",  x"f3",  x"eb",  x"11",  x"00",  x"b7",  x"01",  x"0b", -- 1358
         x"00",  x"ed",  x"b0",  x"af",  x"12",  x"32",  x"96",  x"b7", -- 1360
         x"67",  x"6f",  x"22",  x"97",  x"b7",  x"3e",  x"0d",  x"cd", -- 1368
         x"4a",  x"d1",  x"cb",  x"57",  x"20",  x"40",  x"06",  x"82", -- 1370
         x"21",  x"0c",  x"b7",  x"16",  x"03",  x"1e",  x"0b",  x"ed", -- 1378
         x"78",  x"f5",  x"e6",  x"7f",  x"04",  x"77",  x"23",  x"7b", -- 1380
         x"fe",  x"03",  x"28",  x"01",  x"f1",  x"1d",  x"20",  x"ef", -- 1388
         x"36",  x"00",  x"23",  x"04",  x"f1",  x"77",  x"23",  x"15", -- 1390
         x"20",  x"e3",  x"21",  x"0c",  x"b7",  x"06",  x"03",  x"e5", -- 1398
         x"11",  x"00",  x"b7",  x"1a",  x"a7",  x"c4",  x"28",  x"d4", -- 13A0
         x"e1",  x"d4",  x"d7",  x"d3",  x"11",  x"0d",  x"00",  x"19", -- 13A8
         x"10",  x"ed",  x"3e",  x"05",  x"18",  x"b9",  x"3a",  x"a0", -- 13B0
         x"b7",  x"a7",  x"c4",  x"db",  x"f4",  x"3e",  x"15",  x"cd", -- 13B8
         x"4a",  x"d1",  x"1e",  x"14",  x"06",  x"82",  x"ed",  x"78", -- 13C0
         x"e6",  x"7f",  x"04",  x"f5",  x"cd",  x"d5",  x"f3",  x"f1", -- 13C8
         x"1d",  x"20",  x"f3",  x"2a",  x"97",  x"b7",  x"c9",  x"7e", -- 13D0
         x"fe",  x"20",  x"c8",  x"e5",  x"3a",  x"a0",  x"b7",  x"fe", -- 13D8
         x"27",  x"cc",  x"00",  x"d4",  x"e1",  x"e5",  x"cd",  x"06", -- 13E0
         x"f9",  x"3e",  x"20",  x"cb",  x"7e",  x"28",  x"02",  x"3e", -- 13E8
         x"2a",  x"cd",  x"d5",  x"f3",  x"cd",  x"bc",  x"f3",  x"2a", -- 13F0
         x"97",  x"b7",  x"23",  x"22",  x"97",  x"b7",  x"e1",  x"c9", -- 13F8
         x"21",  x"96",  x"b7",  x"34",  x"3a",  x"9f",  x"b7",  x"3d", -- 1400
         x"96",  x"20",  x"04",  x"77",  x"cd",  x"f6",  x"f3",  x"c3", -- 1408
         x"db",  x"f4",  x"eb",  x"7e",  x"e6",  x"df",  x"cc",  x"67", -- 1410
         x"f5",  x"3f",  x"d0",  x"cd",  x"94",  x"d1",  x"3e",  x"11", -- 1418
         x"cd",  x"4a",  x"d1",  x"d8",  x"18",  x"97",  x"23",  x"13", -- 1420
         x"1a",  x"b6",  x"c8",  x"1a",  x"fe",  x"2a",  x"28",  x"16", -- 1428
         x"fe",  x"01",  x"d8",  x"7e",  x"fe",  x"01",  x"d8",  x"1a", -- 1430
         x"fe",  x"3f",  x"28",  x"ea",  x"cb",  x"6e",  x"cc",  x"3d", -- 1438
         x"f5",  x"be",  x"28",  x"e2",  x"37",  x"c9",  x"e5",  x"d5", -- 1440
         x"cd",  x"27",  x"d4",  x"d1",  x"e1",  x"d0",  x"7e",  x"23", -- 1448
         x"b7",  x"20",  x"f3",  x"37",  x"c9",  x"1a",  x"e6",  x"df", -- 1450
         x"20",  x"13",  x"cd",  x"cf",  x"f0",  x"41",  x"6c",  x"74", -- 1458
         x"65",  x"72",  x"20",  x"00",  x"21",  x"0c",  x"00",  x"cd", -- 1460
         x"a6",  x"d1",  x"d8",  x"18",  x"04",  x"eb",  x"cd",  x"aa", -- 1468
         x"d1",  x"3e",  x"29",  x"cd",  x"4a",  x"d1",  x"d8",  x"1a", -- 1470
         x"e6",  x"df",  x"20",  x"13",  x"cd",  x"cf",  x"f0",  x"4e", -- 1478
         x"65",  x"75",  x"65",  x"72",  x"20",  x"00",  x"21",  x"0c", -- 1480
         x"00",  x"cd",  x"a6",  x"d1",  x"d8",  x"18",  x"04",  x"eb", -- 1488
         x"cd",  x"aa",  x"d1",  x"3e",  x"21",  x"cd",  x"4a",  x"d1", -- 1490
         x"d8",  x"cd",  x"cf",  x"f0",  x"4f",  x"4b",  x"2e",  x"0d", -- 1498
         x"0a",  x"00",  x"c9",  x"7f",  x"7f",  x"54",  x"59",  x"50", -- 14A0
         x"45",  x"1f",  x"cd",  x"c8",  x"d5",  x"d8",  x"cd",  x"c9", -- 14A8
         x"e4",  x"04",  x"38",  x"77",  x"3a",  x"10",  x"b7",  x"fe", -- 14B0
         x"02",  x"38",  x"1b",  x"fe",  x"05",  x"30",  x"17",  x"18", -- 14B8
         x"0f",  x"3e",  x"0c",  x"cd",  x"8c",  x"e0",  x"3e",  x"0a", -- 14C0
         x"cd",  x"8c",  x"e0",  x"7b",  x"fe",  x"80",  x"20",  x"09", -- 14C8
         x"cd",  x"c9",  x"e4",  x"01",  x"38",  x"3f",  x"11",  x"00", -- 14D0
         x"b7",  x"1a",  x"1c",  x"fe",  x"03",  x"28",  x"36",  x"fe", -- 14D8
         x"1a",  x"28",  x"32",  x"fe",  x"20",  x"30",  x"1c",  x"fe", -- 14E0
         x"0a",  x"28",  x"18",  x"fe",  x"0d",  x"28",  x"14",  x"fe", -- 14E8
         x"09",  x"20",  x"0e",  x"3e",  x"20",  x"cd",  x"d5",  x"f3", -- 14F0
         x"3a",  x"a0",  x"b7",  x"e6",  x"07",  x"20",  x"f4",  x"18", -- 14F8
         x"05",  x"3e",  x"2e",  x"cd",  x"d5",  x"f3",  x"3a",  x"a1", -- 1500
         x"b7",  x"3c",  x"21",  x"9f",  x"b7",  x"be",  x"20",  x"bb", -- 1508
         x"cd",  x"e4",  x"d5",  x"20",  x"ac",  x"cd",  x"db",  x"f4", -- 1510
         x"18",  x"11",  x"7f",  x"7f",  x"44",  x"55",  x"4d",  x"50", -- 1518
         x"1f",  x"cd",  x"c8",  x"d5",  x"d8",  x"cd",  x"c9",  x"e4", -- 1520
         x"04",  x"30",  x"25",  x"cd",  x"c9",  x"e4",  x"05",  x"cd", -- 1528
         x"c0",  x"e4",  x"3a",  x"80",  x"b7",  x"32",  x"05",  x"b8", -- 1530
         x"c3",  x"9c",  x"fb",  x"3e",  x"0c",  x"cd",  x"8c",  x"e0", -- 1538
         x"3e",  x"0a",  x"cd",  x"8c",  x"e0",  x"7b",  x"fe",  x"80", -- 1540
         x"20",  x"09",  x"cd",  x"c9",  x"e4",  x"01",  x"38",  x"db", -- 1548
         x"11",  x"00",  x"b7",  x"eb",  x"cd",  x"bc",  x"f3",  x"0e", -- 1550
         x"08",  x"cd",  x"a9",  x"d7",  x"eb",  x"cd",  x"db",  x"f4", -- 1558
         x"3a",  x"a1",  x"b7",  x"3c",  x"21",  x"9f",  x"b7",  x"be", -- 1560
         x"20",  x"db",  x"cd",  x"e4",  x"d5",  x"28",  x"bc",  x"18", -- 1568
         x"ca",  x"49",  x"4e",  x"49",  x"54",  x"49",  x"41",  x"4c", -- 1570
         x"2e",  x"55",  x"55",  x"55",  x"00",  x"7f",  x"7f",  x"49", -- 1578
         x"4e",  x"49",  x"54",  x"1f",  x"1a",  x"e6",  x"df",  x"20", -- 1580
         x"03",  x"11",  x"71",  x"d5",  x"cd",  x"c8",  x"d5",  x"d8", -- 1588
         x"cd",  x"c9",  x"e4",  x"04",  x"38",  x"95",  x"21",  x"00", -- 1590
         x"b7",  x"11",  x"80",  x"a8",  x"7e",  x"a7",  x"28",  x"13", -- 1598
         x"fe",  x"03",  x"28",  x"15",  x"fe",  x"0a",  x"28",  x"0b", -- 15A0
         x"fe",  x"1a",  x"28",  x"0d",  x"12",  x"1c",  x"7b",  x"fe", -- 15A8
         x"7f",  x"28",  x"06",  x"2c",  x"7d",  x"fe",  x"80",  x"20", -- 15B0
         x"e3",  x"af",  x"12",  x"21",  x"80",  x"a8",  x"22",  x"d1", -- 15B8
         x"b7",  x"dd",  x"cb",  x"08",  x"f6",  x"c3",  x"2b",  x"d5", -- 15C0
         x"cd",  x"97",  x"ed",  x"37",  x"c8",  x"eb",  x"7e",  x"e6", -- 15C8
         x"df",  x"cc",  x"67",  x"f5",  x"d8",  x"cd",  x"46",  x"f5", -- 15D0
         x"3a",  x"05",  x"b8",  x"32",  x"80",  x"b7",  x"3e",  x"01", -- 15D8
         x"32",  x"05",  x"b8",  x"c9",  x"cd",  x"f0",  x"f3",  x"fe", -- 15E0
         x"03",  x"c8",  x"fe",  x"0f",  x"c0",  x"cd",  x"d5",  x"f3", -- 15E8
         x"18",  x"f2",  x"fe",  x"08",  x"28",  x"1d",  x"30",  x"26", -- 15F0
         x"4f",  x"87",  x"87",  x"dd",  x"ae",  x"08",  x"e6",  x"1c", -- 15F8
         x"dd",  x"ae",  x"08",  x"47",  x"e6",  x"1c",  x"87",  x"87", -- 1600
         x"87",  x"26",  x"a9",  x"6f",  x"7e",  x"b9",  x"37",  x"c0", -- 1608
         x"dd",  x"70",  x"08",  x"cd",  x"90",  x"ed",  x"f5",  x"21", -- 1610
         x"04",  x"a9",  x"b5",  x"6f",  x"f1",  x"c9",  x"3c",  x"28", -- 1618
         x"0f",  x"cd",  x"13",  x"d6",  x"06",  x"04",  x"7e",  x"23", -- 1620
         x"fe",  x"20",  x"d4",  x"d5",  x"f3",  x"10",  x"f7",  x"c9", -- 1628
         x"21",  x"00",  x"a9",  x"4d",  x"7e",  x"b9",  x"20",  x"12", -- 1630
         x"23",  x"23",  x"23",  x"23",  x"cd",  x"cd",  x"f3",  x"3e", -- 1638
         x"3d",  x"cd",  x"d5",  x"f3",  x"cd",  x"24",  x"d6",  x"cd", -- 1640
         x"db",  x"f4",  x"7d",  x"f6",  x"1f",  x"3c",  x"6f",  x"0c", -- 1648
         x"79",  x"fe",  x"08",  x"20",  x"df",  x"c9",  x"cd",  x"db", -- 1650
         x"f4",  x"cd",  x"30",  x"d6",  x"cd",  x"cf",  x"f0",  x"02", -- 1658
         x"3f",  x"00",  x"cd",  x"f6",  x"f3",  x"fe",  x"30",  x"38", -- 1660
         x"f3",  x"fe",  x"38",  x"30",  x"ef",  x"f5",  x"e6",  x"0f", -- 1668
         x"cd",  x"f2",  x"d5",  x"30",  x"03",  x"f1",  x"18",  x"e4", -- 1670
         x"f1",  x"cd",  x"8c",  x"e0",  x"c3",  x"db",  x"f4",  x"01", -- 1678
         x"f1",  x"83",  x"ed",  x"78",  x"fe",  x"20",  x"30",  x"13", -- 1680
         x"cd",  x"cf",  x"f0",  x"4b",  x"65",  x"69",  x"6e",  x"20", -- 1688
         x"44",  x"45",  x"50",  x"32",  x"21",  x"07",  x"0d",  x"0a", -- 1690
         x"00",  x"37",  x"c9",  x"eb",  x"7e",  x"e6",  x"df",  x"20", -- 1698
         x"2d",  x"cd",  x"cf",  x"f0",  x"44",  x"72",  x"69",  x"76", -- 16A0
         x"65",  x"3a",  x"00",  x"3e",  x"01",  x"cd",  x"83",  x"d1", -- 16A8
         x"01",  x"f1",  x"81",  x"ed",  x"78",  x"cd",  x"d5",  x"f3", -- 16B0
         x"04",  x"ed",  x"78",  x"e6",  x"0f",  x"c4",  x"cd",  x"f3", -- 16B8
         x"3e",  x"06",  x"32",  x"a0",  x"b7",  x"cd",  x"99",  x"f4", -- 16C0
         x"3f",  x"d0",  x"21",  x"06",  x"00",  x"19",  x"01",  x"f1", -- 16C8
         x"81",  x"7e",  x"a7",  x"c8",  x"cd",  x"3d",  x"f5",  x"ed", -- 16D0
         x"79",  x"23",  x"7e",  x"a7",  x"3e",  x"03",  x"28",  x"10", -- 16D8
         x"eb",  x"cd",  x"eb",  x"f4",  x"3e",  x"00",  x"38",  x"03", -- 16E0
         x"3a",  x"97",  x"b7",  x"04",  x"ed",  x"79",  x"3e",  x"07", -- 16E8
         x"cd",  x"83",  x"d1",  x"c9",  x"e6",  x"03",  x"4f",  x"cd", -- 16F0
         x"90",  x"ed",  x"81",  x"81",  x"4f",  x"06",  x"00",  x"21", -- 16F8
         x"18",  x"a9",  x"09",  x"7e",  x"23",  x"66",  x"6f",  x"e9", -- 1700
         x"cd",  x"cf",  x"f0",  x"54",  x"61",  x"70",  x"65",  x"2d", -- 1708
         x"44",  x"69",  x"72",  x"65",  x"63",  x"74",  x"6f",  x"72", -- 1710
         x"79",  x"3a",  x"0d",  x"0a",  x"00",  x"21",  x"00",  x"00", -- 1718
         x"22",  x"97",  x"b7",  x"db",  x"88",  x"f6",  x"60",  x"d3", -- 1720
         x"88",  x"3e",  x"0a",  x"cd",  x"a3",  x"e2",  x"cd",  x"46", -- 1728
         x"f5",  x"dd",  x"36",  x"03",  x"01",  x"cd",  x"c9",  x"e4", -- 1730
         x"01",  x"38",  x"39",  x"dd",  x"7e",  x"02",  x"3d",  x"28", -- 1738
         x"08",  x"cd",  x"c9",  x"f0",  x"2a",  x"19",  x"00",  x"18", -- 1740
         x"2b",  x"cd",  x"3c",  x"f6",  x"2a",  x"97",  x"b7",  x"23", -- 1748
         x"22",  x"97",  x"b7",  x"3a",  x"10",  x"b7",  x"d6",  x"02", -- 1750
         x"fe",  x"08",  x"30",  x"15",  x"2a",  x"11",  x"b7",  x"ed", -- 1758
         x"5b",  x"13",  x"b7",  x"cd",  x"e2",  x"f4",  x"2a",  x"15", -- 1760
         x"b7",  x"3a",  x"10",  x"b7",  x"fe",  x"03",  x"d4",  x"b4", -- 1768
         x"f3",  x"cd",  x"db",  x"f4",  x"cd",  x"7c",  x"e3",  x"30", -- 1770
         x"b8",  x"db",  x"88",  x"e6",  x"9f",  x"d3",  x"88",  x"2a", -- 1778
         x"97",  x"b7",  x"c9",  x"db",  x"88",  x"ee",  x"40",  x"d3", -- 1780
         x"88",  x"c9",  x"e5",  x"d5",  x"e5",  x"23",  x"23",  x"23", -- 1788
         x"11",  x"f5",  x"b7",  x"01",  x"08",  x"00",  x"ed",  x"b0", -- 1790
         x"e1",  x"06",  x"03",  x"7e",  x"23",  x"e6",  x"7f",  x"12", -- 1798
         x"13",  x"10",  x"f8",  x"d1",  x"e1",  x"c9",  x"cd",  x"b4", -- 17A0
         x"f3",  x"e5",  x"41",  x"cd",  x"80",  x"fb",  x"23",  x"cd", -- 17A8
         x"b9",  x"f3",  x"10",  x"f7",  x"e1",  x"41",  x"3e",  x"09", -- 17B0
         x"cd",  x"d5",  x"f3",  x"cd",  x"80",  x"fb",  x"23",  x"cd", -- 17B8
         x"b5",  x"f7",  x"10",  x"f7",  x"c9",  x"0a",  x"0d",  x"09", -- 17C0
         x"1b",  x"4a",  x"18",  x"1b",  x"2a",  x"05",  x"40",  x"01", -- 17C8
         x"0a",  x"0d",  x"09",  x"1b",  x"4a",  x"18",  x"1b",  x"2a", -- 17D0
         x"05",  x"80",  x"02",  x"0e",  x"1b",  x"5b",  x"30",  x"31", -- 17D8
         x"65",  x"1b",  x"5b",  x"31",  x"32",  x"60",  x"1b",  x"4b", -- 17E0
         x"40",  x"01",  x"0e",  x"1b",  x"5b",  x"30",  x"31",  x"65", -- 17E8
         x"1b",  x"5b",  x"31",  x"32",  x"60",  x"1b",  x"4b",  x"80", -- 17F0
         x"02",  x"09",  x"0d",  x"09",  x"1b",  x"4a",  x"18",  x"1b", -- 17F8
         x"4b",  x"40",  x"01",  x"0a",  x"0d",  x"09",  x"1b",  x"4a", -- 1800
         x"18",  x"1b",  x"2a",  x"27",  x"40",  x"01",  x"0a",  x"0d", -- 1808
         x"09",  x"1b",  x"4a",  x"18",  x"1b",  x"2a",  x"00",  x"40", -- 1810
         x"01",  x"0a",  x"0d",  x"09",  x"1b",  x"4a",  x"18",  x"1b", -- 1818
         x"2a",  x"27",  x"c0",  x"03",  x"00",  x"47",  x"5b",  x"04", -- 1820
         x"04",  x"03",  x"20",  x"05",  x"6a",  x"47",  x"2e",  x"18", -- 1828
         x"04",  x"44",  x"03",  x"e1",  x"05",  x"6a",  x"02",  x"0d", -- 1830
         x"02",  x"47",  x"2e",  x"0b",  x"0b",  x"18",  x"02",  x"e2", -- 1838
         x"04",  x"44",  x"03",  x"e1",  x"05",  x"ea",  x"11",  x"18", -- 1840
         x"0b",  x"07",  x"18",  x"04",  x"44",  x"03",  x"e1",  x"05", -- 1848
         x"6a",  x"8c",  x"e0",  x"76",  x"e5",  x"bd",  x"b7",  x"c3", -- 1850
         x"b7",  x"f6",  x"f3",  x"7b",  x"e5",  x"c0",  x"b7",  x"c6", -- 1858
         x"b7",  x"80",  x"e5",  x"85",  x"e5",  x"8a",  x"e5",  x"8f", -- 1860
         x"e5",  x"68",  x"e3",  x"66",  x"f1",  x"73",  x"e3",  x"af", -- 1868
         x"f7",  x"c6",  x"f6",  x"af",  x"f6",  x"69",  x"f2",  x"89", -- 1870
         x"f3",  x"a3",  x"e2",  x"ff",  x"f5",  x"f0",  x"f3",  x"99", -- 1878
         x"f4",  x"eb",  x"f4",  x"d1",  x"f4",  x"b4",  x"f3",  x"e2", -- 1880
         x"f4",  x"c4",  x"f3",  x"5a",  x"f3",  x"8f",  x"f3",  x"9c", -- 1888
         x"f3",  x"8c",  x"f3",  x"99",  x"f3",  x"20",  x"f5",  x"cf", -- 1890
         x"f0",  x"d5",  x"f3",  x"22",  x"f8",  x"04",  x"f1",  x"1d", -- 1898
         x"f1",  x"d4",  x"e2",  x"d6",  x"e2",  x"7c",  x"e3",  x"bc", -- 18A0
         x"f3",  x"db",  x"f4",  x"c0",  x"f3",  x"dd",  x"f7",  x"58", -- 18A8
         x"f8",  x"50",  x"f8",  x"96",  x"fb",  x"68",  x"e0",  x"5c", -- 18B0
         x"e0",  x"4c",  x"e0",  x"0c",  x"f9",  x"85",  x"f5",  x"71", -- 18B8
         x"f8",  x"79",  x"f8",  x"1a",  x"f8",  x"11",  x"f8",  x"cc", -- 18C0
         x"f7",  x"f7",  x"f7",  x"ff",  x"f7",  x"68",  x"f8",  x"60", -- 18C8
         x"f8",  x"8a",  x"ed",  x"ac",  x"fb",  x"b5",  x"f7",  x"4f", -- 18D0
         x"f5",  x"61",  x"f5",  x"06",  x"f9",  x"fc",  x"f1",  x"b9", -- 18D8
         x"f9",  x"e1",  x"f9",  x"d7",  x"fb",  x"ff",  x"05",  x"00", -- 18E0
         x"01",  x"54",  x"41",  x"50",  x"45",  x"0f",  x"d0",  x"72", -- 18E8
         x"d0",  x"00",  x"d0",  x"76",  x"e4",  x"6f",  x"d0",  x"7d", -- 18F0
         x"e4",  x"bf",  x"f4",  x"bf",  x"f4",  x"08",  x"d7",  x"83", -- 18F8
         x"d7",  x"03",  x"f3",  x"03",  x"f3",  x"01",  x"05",  x"00", -- 1900
         x"01",  x"44",  x"49",  x"53",  x"4b",  x"2e",  x"d1",  x"04", -- 1908
         x"d1",  x"24",  x"d1",  x"88",  x"d1",  x"f6",  x"d0",  x"20", -- 1910
         x"d1",  x"bf",  x"f4",  x"bf",  x"f4",  x"5a",  x"d3",  x"7f", -- 1918
         x"d6",  x"12",  x"d4",  x"55",  x"d4",  x"07",  x"8a",  x"01", -- 1920
         x"e4",  x"88",  x"02",  x"1f",  x"0f",  x"8a",  x"02",  x"0f", -- 1928
         x"03",  x"8b",  x"03",  x"e6",  x"0f",  x"83",  x"89",  x"01", -- 1930
         x"ff",  x"84",  x"01",  x"28",  x"86",  x"01",  x"e3",  x"04", -- 1938
         x"8a",  x"01",  x"e4",  x"8b",  x"01",  x"e6",  x"8c",  x"01", -- 1940
         x"e8",  x"8e",  x"02",  x"47",  x"0c",  x"03",  x"06",  x"02", -- 1948
         x"cf",  x"00",  x"07",  x"02",  x"cf",  x"fe",  x"05",  x"01", -- 1950
         x"01",  x"02",  x"0b",  x"0a",  x"0d",  x"08",  x"00",  x"00", -- 1958
         x"0d",  x"09",  x"00",  x"00",  x"20",  x"d5",  x"e3",  x"90", -- 1960
         x"fa",  x"a4",  x"e5",  x"ed",  x"e2",  x"b3",  x"e5",  x"94", -- 1968
         x"e5",  x"ac",  x"ed",  x"e1",  x"e2",  x"7b",  x"7c",  x"7d", -- 1970
         x"7e",  x"5b",  x"5c",  x"5d",  x"84",  x"94",  x"81",  x"e1", -- 1978
         x"8e",  x"99",  x"9a",  x"7f",  x"7f",  x"68",  x"65",  x"6c", -- 1980
         x"70",  x"01",  x"cd",  x"cf",  x"f0",  x"20",  x"4b",  x"43", -- 1988
         x"2d",  x"43",  x"6c",  x"75",  x"62",  x"20",  x"43",  x"41", -- 1990
         x"4f",  x"53",  x"20",  x"34",  x"2e",  x"37",  x"20",  x"31", -- 1998
         x"30",  x"2e",  x"30",  x"34",  x"2e",  x"32",  x"30",  x"31", -- 19A0
         x"39",  x"0d",  x"0a",  x"00",  x"c9",  x"ff",  x"ff",  x"ff", -- 19A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 19B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 19B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 19C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 19C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 19D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 19D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 19E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 19E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 19F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 19F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1A98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1AA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1AA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1AB0
         x"78",  x"60",  x"60",  x"60",  x"60",  x"60",  x"78",  x"00", -- 1AB8
         x"c0",  x"60",  x"30",  x"18",  x"0c",  x"06",  x"02",  x"00", -- 1AC0
         x"78",  x"18",  x"18",  x"18",  x"18",  x"18",  x"78",  x"00", -- 1AC8
         x"30",  x"30",  x"18",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1AD0
         x"1c",  x"30",  x"30",  x"e0",  x"30",  x"30",  x"1c",  x"00", -- 1AD8
         x"18",  x"18",  x"18",  x"00",  x"18",  x"18",  x"18",  x"00", -- 1AE0
         x"e0",  x"30",  x"30",  x"1c",  x"30",  x"30",  x"e0",  x"00", -- 1AE8
         x"76",  x"dc",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1AF0
         x"00",  x"10",  x"38",  x"6c",  x"c6",  x"c6",  x"fe",  x"00", -- 1AF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"81",  x"ff", -- 1B00
         x"7e",  x"81",  x"a5",  x"81",  x"bd",  x"99",  x"81",  x"7e", -- 1B08
         x"7e",  x"ff",  x"db",  x"ff",  x"c3",  x"e7",  x"ff",  x"7e", -- 1B10
         x"6c",  x"fe",  x"fe",  x"fe",  x"7c",  x"38",  x"10",  x"00", -- 1B18
         x"10",  x"38",  x"7c",  x"fe",  x"7c",  x"38",  x"10",  x"00", -- 1B20
         x"38",  x"7c",  x"38",  x"fe",  x"fe",  x"7c",  x"38",  x"7c", -- 1B28
         x"10",  x"10",  x"38",  x"7c",  x"fe",  x"7c",  x"38",  x"7c", -- 1B30
         x"00",  x"00",  x"18",  x"3c",  x"3c",  x"18",  x"00",  x"00", -- 1B38
         x"ff",  x"ff",  x"e7",  x"c3",  x"c3",  x"e7",  x"ff",  x"ff", -- 1B40
         x"00",  x"3c",  x"66",  x"42",  x"42",  x"66",  x"3c",  x"00", -- 1B48
         x"ff",  x"c3",  x"99",  x"bd",  x"bd",  x"99",  x"c3",  x"ff", -- 1B50
         x"0f",  x"07",  x"0f",  x"7d",  x"cc",  x"cc",  x"cc",  x"78", -- 1B58
         x"3c",  x"66",  x"66",  x"66",  x"3c",  x"18",  x"7e",  x"18", -- 1B60
         x"3f",  x"33",  x"3f",  x"30",  x"30",  x"70",  x"f0",  x"e0", -- 1B68
         x"7f",  x"63",  x"7f",  x"63",  x"63",  x"67",  x"e6",  x"c0", -- 1B70
         x"99",  x"5a",  x"3c",  x"e7",  x"e7",  x"3c",  x"5a",  x"99", -- 1B78
         x"80",  x"e0",  x"f8",  x"fe",  x"f8",  x"e0",  x"80",  x"00", -- 1B80
         x"02",  x"0e",  x"3e",  x"fe",  x"3e",  x"0e",  x"02",  x"00", -- 1B88
         x"18",  x"3c",  x"7e",  x"18",  x"18",  x"7e",  x"3c",  x"18", -- 1B90
         x"66",  x"66",  x"66",  x"66",  x"66",  x"00",  x"66",  x"00", -- 1B98
         x"7b",  x"db",  x"db",  x"7b",  x"1b",  x"1b",  x"1b",  x"00", -- 1BA0
         x"3c",  x"66",  x"38",  x"6c",  x"6c",  x"38",  x"cc",  x"78", -- 1BA8
         x"00",  x"00",  x"00",  x"00",  x"7e",  x"7e",  x"7e",  x"00", -- 1BB0
         x"18",  x"3c",  x"7e",  x"18",  x"7e",  x"3c",  x"18",  x"ff", -- 1BB8
         x"18",  x"3c",  x"7e",  x"18",  x"18",  x"18",  x"18",  x"00", -- 1BC0
         x"18",  x"18",  x"18",  x"18",  x"7e",  x"3c",  x"18",  x"00", -- 1BC8
         x"00",  x"08",  x"0c",  x"fe",  x"fe",  x"0c",  x"08",  x"00", -- 1BD0
         x"00",  x"20",  x"60",  x"fe",  x"fe",  x"60",  x"20",  x"00", -- 1BD8
         x"00",  x"00",  x"c0",  x"c0",  x"c0",  x"fe",  x"00",  x"00", -- 1BE0
         x"00",  x"24",  x"66",  x"ff",  x"ff",  x"66",  x"24",  x"00", -- 1BE8
         x"00",  x"18",  x"3c",  x"7e",  x"ff",  x"ff",  x"00",  x"00", -- 1BF0
         x"00",  x"ff",  x"ff",  x"7e",  x"3c",  x"18",  x"00",  x"00", -- 1BF8
         x"78",  x"cc",  x"c0",  x"c0",  x"cc",  x"78",  x"10",  x"70", -- 1C00
         x"00",  x"cc",  x"00",  x"cc",  x"cc",  x"cc",  x"76",  x"00", -- 1C08
         x"1c",  x"00",  x"78",  x"cc",  x"fc",  x"c0",  x"78",  x"00", -- 1C10
         x"78",  x"84",  x"78",  x"0c",  x"7c",  x"cc",  x"76",  x"00", -- 1C18
         x"6c",  x"00",  x"78",  x"0c",  x"7c",  x"cc",  x"76",  x"00", -- 1C20
         x"e0",  x"00",  x"78",  x"0c",  x"7c",  x"cc",  x"76",  x"00", -- 1C28
         x"30",  x"30",  x"78",  x"0c",  x"7c",  x"cc",  x"76",  x"00", -- 1C30
         x"00",  x"78",  x"cc",  x"c0",  x"cc",  x"78",  x"10",  x"70", -- 1C38
         x"78",  x"84",  x"78",  x"cc",  x"fc",  x"c0",  x"78",  x"00", -- 1C40
         x"cc",  x"00",  x"78",  x"cc",  x"fc",  x"c0",  x"78",  x"00", -- 1C48
         x"e0",  x"00",  x"78",  x"cc",  x"fc",  x"c0",  x"78",  x"00", -- 1C50
         x"d8",  x"00",  x"70",  x"30",  x"30",  x"30",  x"78",  x"00", -- 1C58
         x"70",  x"88",  x"70",  x"30",  x"30",  x"30",  x"78",  x"00", -- 1C60
         x"e0",  x"00",  x"70",  x"30",  x"30",  x"30",  x"78",  x"00", -- 1C68
         x"cc",  x"30",  x"78",  x"cc",  x"fc",  x"cc",  x"cc",  x"00", -- 1C70
         x"78",  x"84",  x"30",  x"78",  x"cc",  x"fc",  x"cc",  x"00", -- 1C78
         x"1c",  x"00",  x"fc",  x"60",  x"78",  x"60",  x"fc",  x"00", -- 1C80
         x"00",  x"00",  x"6c",  x"92",  x"9e",  x"90",  x"7e",  x"00", -- 1C88
         x"3e",  x"78",  x"d8",  x"fe",  x"d8",  x"d8",  x"de",  x"00", -- 1C90
         x"78",  x"84",  x"00",  x"78",  x"cc",  x"cc",  x"78",  x"00", -- 1C98
         x"00",  x"cc",  x"00",  x"78",  x"cc",  x"cc",  x"78",  x"00", -- 1CA0
         x"00",  x"e0",  x"00",  x"78",  x"cc",  x"cc",  x"78",  x"00", -- 1CA8
         x"78",  x"84",  x"00",  x"cc",  x"cc",  x"cc",  x"76",  x"00", -- 1CB0
         x"00",  x"e0",  x"00",  x"cc",  x"cc",  x"cc",  x"76",  x"00", -- 1CB8
         x"00",  x"cc",  x"00",  x"cc",  x"cc",  x"7c",  x"0c",  x"f8", -- 1CC0
         x"c6",  x"38",  x"6c",  x"c6",  x"c6",  x"6c",  x"38",  x"00", -- 1CC8
         x"cc",  x"00",  x"cc",  x"cc",  x"cc",  x"cc",  x"78",  x"00", -- 1CD0
         x"00",  x"10",  x"7c",  x"d6",  x"d0",  x"d6",  x"7c",  x"10", -- 1CD8
         x"38",  x"6c",  x"64",  x"f0",  x"60",  x"e6",  x"fc",  x"00", -- 1CE0
         x"66",  x"66",  x"3c",  x"7e",  x"18",  x"7e",  x"18",  x"18", -- 1CE8
         x"f8",  x"cc",  x"cc",  x"fa",  x"c6",  x"cf",  x"c6",  x"c7", -- 1CF0
         x"0e",  x"1b",  x"18",  x"3c",  x"18",  x"18",  x"d8",  x"70", -- 1CF8
         x"1c",  x"00",  x"78",  x"0c",  x"7c",  x"cc",  x"76",  x"00", -- 1D00
         x"38",  x"00",  x"70",  x"30",  x"30",  x"30",  x"78",  x"00", -- 1D08
         x"00",  x"1c",  x"00",  x"78",  x"cc",  x"cc",  x"78",  x"00", -- 1D10
         x"00",  x"1c",  x"00",  x"cc",  x"cc",  x"cc",  x"76",  x"00", -- 1D18
         x"00",  x"f8",  x"00",  x"f8",  x"cc",  x"cc",  x"cc",  x"00", -- 1D20
         x"fc",  x"00",  x"cc",  x"ec",  x"fc",  x"dc",  x"cc",  x"00", -- 1D28
         x"00",  x"3c",  x"6c",  x"6c",  x"3e",  x"00",  x"7e",  x"00", -- 1D30
         x"00",  x"38",  x"6c",  x"6c",  x"38",  x"00",  x"7c",  x"00", -- 1D38
         x"30",  x"00",  x"30",  x"18",  x"0c",  x"cc",  x"78",  x"00", -- 1D40
         x"00",  x"00",  x"00",  x"7e",  x"60",  x"60",  x"00",  x"00", -- 1D48
         x"00",  x"00",  x"00",  x"7e",  x"06",  x"06",  x"00",  x"00", -- 1D50
         x"c3",  x"c6",  x"cc",  x"de",  x"33",  x"66",  x"cc",  x"0f", -- 1D58
         x"c3",  x"c6",  x"cc",  x"db",  x"37",  x"6f",  x"cf",  x"03", -- 1D60
         x"30",  x"00",  x"30",  x"30",  x"78",  x"78",  x"30",  x"00", -- 1D68
         x"00",  x"33",  x"66",  x"cc",  x"66",  x"33",  x"00",  x"00", -- 1D70
         x"00",  x"cc",  x"66",  x"33",  x"66",  x"cc",  x"00",  x"00", -- 1D78
         x"22",  x"88",  x"22",  x"88",  x"22",  x"88",  x"22",  x"88", -- 1D80
         x"55",  x"aa",  x"55",  x"aa",  x"55",  x"aa",  x"55",  x"aa", -- 1D88
         x"77",  x"dd",  x"77",  x"dd",  x"77",  x"dd",  x"77",  x"dd", -- 1D90
         x"18",  x"18",  x"18",  x"18",  x"18",  x"18",  x"18",  x"18", -- 1D98
         x"18",  x"18",  x"18",  x"f8",  x"18",  x"18",  x"18",  x"18", -- 1DA0
         x"18",  x"18",  x"f8",  x"18",  x"f8",  x"18",  x"18",  x"18", -- 1DA8
         x"36",  x"36",  x"36",  x"f6",  x"36",  x"36",  x"36",  x"36", -- 1DB0
         x"00",  x"00",  x"00",  x"fe",  x"36",  x"36",  x"36",  x"36", -- 1DB8
         x"00",  x"00",  x"f8",  x"18",  x"f8",  x"18",  x"18",  x"18", -- 1DC0
         x"36",  x"36",  x"f6",  x"06",  x"f6",  x"36",  x"36",  x"36", -- 1DC8
         x"36",  x"36",  x"36",  x"36",  x"36",  x"36",  x"36",  x"36", -- 1DD0
         x"00",  x"00",  x"fe",  x"06",  x"f6",  x"36",  x"36",  x"36", -- 1DD8
         x"36",  x"36",  x"f6",  x"06",  x"fe",  x"00",  x"00",  x"00", -- 1DE0
         x"36",  x"36",  x"36",  x"fe",  x"00",  x"00",  x"00",  x"00", -- 1DE8
         x"18",  x"18",  x"f8",  x"18",  x"f8",  x"00",  x"00",  x"00", -- 1DF0
         x"00",  x"00",  x"00",  x"f8",  x"18",  x"18",  x"18",  x"18", -- 1DF8
         x"18",  x"18",  x"18",  x"1f",  x"00",  x"00",  x"00",  x"00", -- 1E00
         x"18",  x"18",  x"18",  x"ff",  x"00",  x"00",  x"00",  x"00", -- 1E08
         x"00",  x"00",  x"00",  x"ff",  x"18",  x"18",  x"18",  x"18", -- 1E10
         x"18",  x"18",  x"18",  x"1f",  x"18",  x"18",  x"18",  x"18", -- 1E18
         x"00",  x"00",  x"00",  x"ff",  x"00",  x"00",  x"00",  x"00", -- 1E20
         x"18",  x"18",  x"18",  x"ff",  x"18",  x"18",  x"18",  x"18", -- 1E28
         x"18",  x"18",  x"1f",  x"18",  x"1f",  x"18",  x"18",  x"18", -- 1E30
         x"36",  x"36",  x"36",  x"37",  x"36",  x"36",  x"36",  x"36", -- 1E38
         x"36",  x"36",  x"37",  x"30",  x"3f",  x"00",  x"00",  x"00", -- 1E40
         x"00",  x"00",  x"3f",  x"30",  x"37",  x"36",  x"36",  x"36", -- 1E48
         x"36",  x"36",  x"f7",  x"00",  x"ff",  x"00",  x"00",  x"00", -- 1E50
         x"00",  x"00",  x"ff",  x"00",  x"f7",  x"36",  x"36",  x"36", -- 1E58
         x"36",  x"36",  x"37",  x"30",  x"37",  x"36",  x"36",  x"36", -- 1E60
         x"00",  x"00",  x"ff",  x"00",  x"ff",  x"00",  x"00",  x"00", -- 1E68
         x"36",  x"36",  x"f7",  x"00",  x"f7",  x"36",  x"36",  x"36", -- 1E70
         x"18",  x"18",  x"ff",  x"00",  x"ff",  x"00",  x"00",  x"00", -- 1E78
         x"36",  x"36",  x"36",  x"ff",  x"00",  x"00",  x"00",  x"00", -- 1E80
         x"00",  x"00",  x"ff",  x"00",  x"ff",  x"18",  x"18",  x"18", -- 1E88
         x"00",  x"00",  x"00",  x"ff",  x"36",  x"36",  x"36",  x"36", -- 1E90
         x"36",  x"36",  x"36",  x"3f",  x"00",  x"00",  x"00",  x"00", -- 1E98
         x"18",  x"18",  x"1f",  x"18",  x"1f",  x"00",  x"00",  x"00", -- 1EA0
         x"00",  x"00",  x"1f",  x"18",  x"1f",  x"18",  x"18",  x"18", -- 1EA8
         x"00",  x"00",  x"00",  x"3f",  x"36",  x"36",  x"36",  x"36", -- 1EB0
         x"36",  x"36",  x"36",  x"ff",  x"36",  x"36",  x"36",  x"36", -- 1EB8
         x"18",  x"18",  x"ff",  x"18",  x"ff",  x"18",  x"18",  x"18", -- 1EC0
         x"18",  x"18",  x"18",  x"f8",  x"00",  x"00",  x"00",  x"00", -- 1EC8
         x"00",  x"00",  x"00",  x"1f",  x"18",  x"18",  x"18",  x"18", -- 1ED0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1ED8
         x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"ff",  x"ff", -- 1EE0
         x"f0",  x"f0",  x"f0",  x"f0",  x"f0",  x"f0",  x"f0",  x"f0", -- 1EE8
         x"0f",  x"0f",  x"0f",  x"0f",  x"0f",  x"0f",  x"0f",  x"0f", -- 1EF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"00",  x"00",  x"00",  x"00", -- 1EF8
         x"00",  x"00",  x"76",  x"dc",  x"cc",  x"dc",  x"76",  x"00", -- 1F00
         x"3c",  x"66",  x"66",  x"6c",  x"66",  x"66",  x"6c",  x"f0", -- 1F08
         x"fe",  x"62",  x"60",  x"60",  x"60",  x"60",  x"f0",  x"00", -- 1F10
         x"00",  x"fe",  x"6c",  x"6c",  x"6c",  x"6c",  x"6e",  x"00", -- 1F18
         x"fc",  x"c4",  x"60",  x"30",  x"60",  x"c4",  x"fc",  x"00", -- 1F20
         x"00",  x"00",  x"7e",  x"d8",  x"d8",  x"d8",  x"70",  x"00", -- 1F28
         x"00",  x"00",  x"cc",  x"cc",  x"cc",  x"f6",  x"c0",  x"c0", -- 1F30
         x"00",  x"7e",  x"d8",  x"18",  x"18",  x"18",  x"18",  x"00", -- 1F38
         x"78",  x"30",  x"78",  x"cc",  x"cc",  x"78",  x"30",  x"78", -- 1F40
         x"38",  x"6c",  x"c6",  x"fe",  x"c6",  x"6c",  x"38",  x"00", -- 1F48
         x"38",  x"6c",  x"c6",  x"c6",  x"6c",  x"6c",  x"ee",  x"00", -- 1F50
         x"1c",  x"30",  x"18",  x"7c",  x"cc",  x"cc",  x"78",  x"00", -- 1F58
         x"00",  x"6c",  x"fe",  x"92",  x"fe",  x"6c",  x"00",  x"00", -- 1F60
         x"03",  x"7e",  x"cc",  x"de",  x"f6",  x"66",  x"fc",  x"80", -- 1F68
         x"3c",  x"60",  x"c0",  x"fc",  x"c0",  x"60",  x"3c",  x"00", -- 1F70
         x"78",  x"cc",  x"cc",  x"cc",  x"cc",  x"cc",  x"cc",  x"00", -- 1F78
         x"00",  x"7e",  x"00",  x"7e",  x"00",  x"7e",  x"00",  x"00", -- 1F80
         x"18",  x"18",  x"7e",  x"18",  x"18",  x"00",  x"7e",  x"00", -- 1F88
         x"30",  x"18",  x"0c",  x"18",  x"30",  x"00",  x"7e",  x"00", -- 1F90
         x"0c",  x"18",  x"30",  x"18",  x"0c",  x"00",  x"7e",  x"00", -- 1F98
         x"0e",  x"1b",  x"1b",  x"18",  x"18",  x"18",  x"18",  x"18", -- 1FA0
         x"18",  x"18",  x"18",  x"18",  x"18",  x"d8",  x"d8",  x"70", -- 1FA8
         x"18",  x"18",  x"00",  x"7e",  x"00",  x"18",  x"18",  x"00", -- 1FB0
         x"00",  x"76",  x"dc",  x"00",  x"76",  x"dc",  x"00",  x"00", -- 1FB8
         x"38",  x"6c",  x"6c",  x"38",  x"00",  x"00",  x"00",  x"00", -- 1FC0
         x"00",  x"00",  x"00",  x"18",  x"18",  x"00",  x"00",  x"00", -- 1FC8
         x"00",  x"00",  x"00",  x"00",  x"18",  x"00",  x"00",  x"00", -- 1FD0
         x"0f",  x"0c",  x"0c",  x"0c",  x"cc",  x"6c",  x"3c",  x"1c", -- 1FD8
         x"78",  x"6c",  x"6c",  x"6c",  x"6c",  x"00",  x"00",  x"00", -- 1FE0
         x"70",  x"18",  x"30",  x"60",  x"78",  x"00",  x"00",  x"00", -- 1FE8
         x"00",  x"00",  x"3c",  x"3c",  x"3c",  x"3c",  x"00",  x"00", -- 1FF0
         x"ff",  x"81",  x"81",  x"81",  x"81",  x"81",  x"81",  x"ff"  -- 1FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
