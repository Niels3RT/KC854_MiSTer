library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_m027 is
    generic(
        ADDR_WIDTH   : integer := 13
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom_m027;

architecture rtl of rom_m027 is
    type rom8192x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom8192x8 := (
         x"7f",  x"7f",  x"45",  x"44",  x"41",  x"53",  x"01",  x"21", -- 0000
         x"00",  x"02",  x"23",  x"cb",  x"7c",  x"20",  x"08",  x"7e", -- 0008
         x"2f",  x"77",  x"be",  x"2f",  x"77",  x"28",  x"f3",  x"2b", -- 0010
         x"e5",  x"cd",  x"03",  x"f0",  x"23",  x"12",  x"0c",  x"0a", -- 0018
         x"0a",  x"3e",  x"3e",  x"3e",  x"20",  x"4b",  x"43",  x"2d", -- 0020
         x"45",  x"44",  x"49",  x"54",  x"4f",  x"52",  x"2f",  x"41", -- 0028
         x"53",  x"53",  x"45",  x"4d",  x"42",  x"4c",  x"45",  x"52", -- 0030
         x"20",  x"3c",  x"3c",  x"3c",  x"0d",  x"0a",  x"0a",  x"4d", -- 0038
         x"45",  x"4d",  x"4f",  x"52",  x"59",  x"20",  x"45",  x"4e", -- 0040
         x"44",  x"20",  x"3a",  x"00",  x"cd",  x"03",  x"f0",  x"1a", -- 0048
         x"01",  x"0f",  x"0c",  x"78",  x"32",  x"a0",  x"b7",  x"cd", -- 0050
         x"7a",  x"c5",  x"eb",  x"cd",  x"03",  x"f0",  x"18",  x"e1", -- 0058
         x"38",  x"b6",  x"e5",  x"ed",  x"5b",  x"97",  x"b7",  x"ed", -- 0060
         x"52",  x"e1",  x"38",  x"ac",  x"eb",  x"23",  x"22",  x"72", -- 0068
         x"00",  x"cb",  x"3c",  x"7c",  x"cb",  x"3c",  x"84",  x"67", -- 0070
         x"2e",  x"00",  x"22",  x"70",  x"00",  x"01",  x"00",  x"02", -- 0078
         x"37",  x"ed",  x"42",  x"eb",  x"38",  x"92",  x"2a",  x"70", -- 0080
         x"00",  x"2b",  x"36",  x"03",  x"22",  x"42",  x"00",  x"22", -- 0088
         x"46",  x"00",  x"60",  x"69",  x"22",  x"40",  x"00",  x"22", -- 0090
         x"44",  x"00",  x"af",  x"67",  x"6f",  x"32",  x"4a",  x"00", -- 0098
         x"22",  x"6e",  x"00",  x"22",  x"48",  x"00",  x"21",  x"00", -- 00A0
         x"b9",  x"1e",  x"03",  x"01",  x"80",  x"00",  x"ed",  x"b1", -- 00A8
         x"e2",  x"b6",  x"c0",  x"1d",  x"20",  x"f8",  x"11",  x"03", -- 00B0
         x"b9",  x"01",  x"7c",  x"00",  x"ed",  x"b0",  x"21",  x"7d", -- 00B8
         x"b9",  x"01",  x"7c",  x"00",  x"ed",  x"b8",  x"36",  x"05", -- 00C0
         x"23",  x"77",  x"23",  x"36",  x"06",  x"23",  x"77",  x"18", -- 00C8
         x"09",  x"7f",  x"7f",  x"52",  x"45",  x"45",  x"44",  x"41", -- 00D0
         x"53",  x"01",  x"dd",  x"36",  x"09",  x"dd",  x"cd",  x"9f", -- 00D8
         x"c1",  x"cd",  x"03",  x"f0",  x"23",  x"0c",  x"0a",  x"3e", -- 00E0
         x"3e",  x"3e",  x"20",  x"45",  x"44",  x"41",  x"53",  x"20", -- 00E8
         x"56",  x"31",  x"2e",  x"34",  x"20",  x"3c",  x"3c",  x"3c", -- 00F0
         x"20",  x"20",  x"20",  x"20",  x"20",  x"46",  x"52",  x"45", -- 00F8
         x"45",  x"20",  x"3a",  x"0d",  x"0a",  x"00",  x"06",  x"28", -- 0100
         x"cd",  x"03",  x"f0",  x"23",  x"5f",  x"00",  x"10",  x"f8", -- 0108
         x"18",  x"0e",  x"dd",  x"dd",  x"4d",  x"45",  x"4e",  x"55", -- 0110
         x"01",  x"e1",  x"cd",  x"03",  x"f0",  x"23",  x"0c",  x"00", -- 0118
         x"cd",  x"b6",  x"c1",  x"cd",  x"03",  x"f0",  x"2d",  x"21", -- 0120
         x"00",  x"ba",  x"01",  x"00",  x"26",  x"cd",  x"03",  x"f0", -- 0128
         x"23",  x"2a",  x"00",  x"cd",  x"03",  x"f0",  x"2a",  x"38", -- 0130
         x"31",  x"dd",  x"7e",  x"09",  x"ed",  x"b1",  x"e2",  x"6a", -- 0138
         x"c1",  x"ed",  x"a1",  x"20",  x"f7",  x"7e",  x"fe",  x"02", -- 0140
         x"38",  x"10",  x"fe",  x"30",  x"38",  x"0c",  x"fe",  x"5f", -- 0148
         x"30",  x"08",  x"cd",  x"03",  x"f0",  x"24",  x"23",  x"0b", -- 0150
         x"18",  x"eb",  x"cd",  x"03",  x"f0",  x"2c",  x"18",  x"cd", -- 0158
         x"cd",  x"b6",  x"c1",  x"cd",  x"03",  x"f0",  x"23",  x"0d", -- 0160
         x"2a",  x"00",  x"cd",  x"03",  x"f0",  x"17",  x"13",  x"1a", -- 0168
         x"fe",  x"20",  x"28",  x"ef",  x"a7",  x"28",  x"ec",  x"dd", -- 0170
         x"7e",  x"09",  x"21",  x"00",  x"ba",  x"01",  x"00",  x"26", -- 0178
         x"cd",  x"03",  x"f0",  x"1d",  x"30",  x"08",  x"e5",  x"cd", -- 0180
         x"03",  x"f0",  x"22",  x"30",  x"07",  x"e1",  x"cd",  x"03", -- 0188
         x"f0",  x"19",  x"18",  x"cf",  x"21",  x"60",  x"c1",  x"e3", -- 0190
         x"23",  x"e5",  x"cd",  x"03",  x"f0",  x"15",  x"c9",  x"21", -- 0198
         x"00",  x"01",  x"22",  x"9c",  x"b7",  x"21",  x"28",  x"1e", -- 01A0
         x"22",  x"9e",  x"b7",  x"cd",  x"03",  x"f0",  x"20",  x"cd", -- 01A8
         x"03",  x"f0",  x"23",  x"12",  x"00",  x"c9",  x"2a",  x"a0", -- 01B0
         x"b7",  x"e5",  x"cd",  x"9f",  x"c1",  x"21",  x"1c",  x"01", -- 01B8
         x"22",  x"a0",  x"b7",  x"ed",  x"5b",  x"44",  x"00",  x"2a", -- 01C0
         x"46",  x"00",  x"af",  x"ed",  x"52",  x"cd",  x"03",  x"f0", -- 01C8
         x"1a",  x"3e",  x"05",  x"32",  x"9d",  x"b7",  x"3e",  x"1a", -- 01D0
         x"32",  x"9f",  x"b7",  x"e1",  x"22",  x"a0",  x"b7",  x"c9", -- 01D8
         x"dd",  x"dd",  x"45",  x"58",  x"49",  x"54",  x"01",  x"3e", -- 01E0
         x"01",  x"32",  x"9d",  x"b7",  x"3e",  x"1e",  x"32",  x"9f", -- 01E8
         x"b7",  x"3a",  x"a1",  x"b7",  x"c6",  x"04",  x"32",  x"a1", -- 01F0
         x"b7",  x"dd",  x"36",  x"09",  x"7f",  x"e1",  x"c9",  x"dd", -- 01F8
         x"dd",  x"43",  x"4c",  x"45",  x"41",  x"52",  x"01",  x"cd", -- 0200
         x"03",  x"f0",  x"23",  x"0d",  x"44",  x"45",  x"4c",  x"45", -- 0208
         x"54",  x"45",  x"20",  x"41",  x"4c",  x"4c",  x"00",  x"cd", -- 0210
         x"56",  x"c5",  x"d8",  x"2a",  x"40",  x"00",  x"22",  x"44", -- 0218
         x"00",  x"2a",  x"42",  x"00",  x"22",  x"46",  x"00",  x"11", -- 0220
         x"00",  x"00",  x"ed",  x"53",  x"48",  x"00",  x"c9",  x"dd", -- 0228
         x"dd",  x"53",  x"41",  x"56",  x"45",  x"01",  x"cd",  x"27", -- 0230
         x"c2",  x"cd",  x"c2",  x"c7",  x"cd",  x"fe",  x"c5",  x"ed", -- 0238
         x"5b",  x"46",  x"00",  x"2a",  x"42",  x"00",  x"af",  x"ed", -- 0240
         x"52",  x"c8",  x"e5",  x"cd",  x"e6",  x"c5",  x"d1",  x"38", -- 0248
         x"46",  x"d5",  x"11",  x"00",  x"b7",  x"dd",  x"73",  x"05", -- 0250
         x"dd",  x"72",  x"06",  x"01",  x"0b",  x"00",  x"ed",  x"b0", -- 0258
         x"cd",  x"03",  x"f0",  x"08",  x"2a",  x"46",  x"00",  x"dd", -- 0260
         x"75",  x"05",  x"dd",  x"74",  x"06",  x"dd",  x"7e",  x"02", -- 0268
         x"cd",  x"03",  x"f0",  x"1c",  x"cd",  x"03",  x"f0",  x"23", -- 0270
         x"20",  x"20",  x"00",  x"e1",  x"01",  x"a0",  x"00",  x"cd", -- 0278
         x"03",  x"f0",  x"2a",  x"38",  x"0e",  x"11",  x"80",  x"00", -- 0280
         x"ed",  x"52",  x"38",  x"07",  x"e5",  x"cd",  x"03",  x"f0", -- 0288
         x"01",  x"18",  x"d4",  x"cd",  x"03",  x"f0",  x"09",  x"cd", -- 0290
         x"03",  x"f0",  x"2c",  x"c9",  x"dd",  x"dd",  x"4c",  x"4f", -- 0298
         x"41",  x"44",  x"01",  x"cd",  x"e6",  x"c5",  x"38",  x"ef", -- 02A0
         x"cd",  x"27",  x"c2",  x"e5",  x"21",  x"00",  x"b7",  x"dd", -- 02A8
         x"75",  x"05",  x"dd",  x"74",  x"06",  x"cd",  x"03",  x"f0", -- 02B0
         x"0a",  x"af",  x"3e",  x"01",  x"cd",  x"49",  x"c3",  x"38", -- 02B8
         x"74",  x"e1",  x"e5",  x"11",  x"00",  x"b7",  x"01",  x"01", -- 02C0
         x"0b",  x"1a",  x"b7",  x"20",  x"02",  x"3e",  x"20",  x"be", -- 02C8
         x"28",  x"07",  x"86",  x"fe",  x"20",  x"28",  x"02",  x"96", -- 02D0
         x"0c",  x"13",  x"23",  x"cd",  x"03",  x"f0",  x"24",  x"10", -- 02D8
         x"e8",  x"cd",  x"03",  x"f0",  x"2c",  x"0d",  x"20",  x"d2", -- 02E0
         x"3e",  x"02",  x"ed",  x"5b",  x"44",  x"00",  x"2a",  x"46", -- 02E8
         x"00",  x"a7",  x"ed",  x"52",  x"28",  x"4d",  x"e5",  x"cd", -- 02F0
         x"49",  x"c3",  x"e1",  x"38",  x"28",  x"01",  x"80",  x"00", -- 02F8
         x"ed",  x"42",  x"30",  x"03",  x"09",  x"44",  x"4d",  x"cd", -- 0300
         x"03",  x"f0",  x"1c",  x"cd",  x"03",  x"f0",  x"23",  x"3e", -- 0308
         x"20",  x"00",  x"21",  x"00",  x"b7",  x"3e",  x"03",  x"be", -- 0310
         x"28",  x"0b",  x"ed",  x"a0",  x"ea",  x"17",  x"c3",  x"dd", -- 0318
         x"7e",  x"02",  x"3c",  x"20",  x"c9",  x"2a",  x"44",  x"00", -- 0320
         x"eb",  x"cd",  x"ea",  x"c7",  x"2a",  x"42",  x"00",  x"2b", -- 0328
         x"36",  x"0a",  x"2b",  x"36",  x"0d",  x"e1",  x"cd",  x"03", -- 0330
         x"f0",  x"0b",  x"3a",  x"4a",  x"00",  x"b7",  x"c8",  x"cd", -- 0338
         x"6a",  x"c7",  x"c9",  x"3c",  x"32",  x"4a",  x"00",  x"18", -- 0340
         x"dc",  x"67",  x"28",  x"09",  x"cd",  x"03",  x"f0",  x"2a", -- 0348
         x"d8",  x"cd",  x"03",  x"f0",  x"05",  x"dd",  x"7e",  x"02", -- 0350
         x"30",  x"15",  x"cd",  x"03",  x"f0",  x"1c",  x"cd",  x"03", -- 0358
         x"f0",  x"23",  x"2a",  x"20",  x"00",  x"7c",  x"3d",  x"20", -- 0360
         x"e3",  x"cd",  x"03",  x"f0",  x"2c",  x"18",  x"dd",  x"bc", -- 0368
         x"c8",  x"fe",  x"ff",  x"20",  x"e5",  x"6c",  x"2d",  x"28", -- 0370
         x"e1",  x"c9",  x"dd",  x"dd",  x"50",  x"52",  x"49",  x"4e", -- 0378
         x"54",  x"01",  x"01",  x"00",  x"01",  x"3a",  x"81",  x"b7", -- 0380
         x"b7",  x"28",  x"0c",  x"45",  x"3d",  x"28",  x"08",  x"4b", -- 0388
         x"21",  x"00",  x"c4",  x"cd",  x"03",  x"f0",  x"1e",  x"c5", -- 0390
         x"cd",  x"27",  x"c2",  x"cd",  x"c2",  x"c7",  x"c1",  x"c5", -- 0398
         x"2a",  x"46",  x"00",  x"16",  x"00",  x"2b",  x"23",  x"7e", -- 03A0
         x"23",  x"fe",  x"03",  x"28",  x"11",  x"fe",  x"0d",  x"28", -- 03A8
         x"16",  x"1e",  x"00",  x"c5",  x"cd",  x"ef",  x"d1",  x"c1", -- 03B0
         x"cd",  x"03",  x"f0",  x"2a",  x"30",  x"e9",  x"cd",  x"03", -- 03B8
         x"f0",  x"23",  x"0d",  x"0a",  x"00",  x"c1",  x"c9",  x"10", -- 03C0
         x"dd",  x"cd",  x"ef",  x"d1",  x"e3",  x"79",  x"b7",  x"28", -- 03C8
         x"2b",  x"0d",  x"20",  x"28",  x"3e",  x"0c",  x"cd",  x"ef", -- 03D0
         x"d1",  x"e5",  x"cd",  x"03",  x"f0",  x"20",  x"cd",  x"03", -- 03D8
         x"f0",  x"23",  x"4e",  x"45",  x"58",  x"54",  x"20",  x"50", -- 03E0
         x"41",  x"47",  x"45",  x"00",  x"cd",  x"56",  x"c5",  x"e1", -- 03E8
         x"38",  x"d3",  x"e5",  x"21",  x"00",  x"c4",  x"cd",  x"03", -- 03F0
         x"f0",  x"1e",  x"e1",  x"4d",  x"44",  x"e3",  x"18",  x"a7", -- 03F8
         x"02",  x"dd",  x"dd",  x"41",  x"53",  x"4d",  x"01",  x"cd", -- 0400
         x"27",  x"c2",  x"cd",  x"c2",  x"c7",  x"af",  x"32",  x"6d", -- 0408
         x"00",  x"cd",  x"03",  x"f0",  x"23",  x"4f",  x"50",  x"54", -- 0410
         x"49",  x"4f",  x"4e",  x"53",  x"28",  x"2b",  x"2c",  x"32", -- 0418
         x"2c",  x"42",  x"2c",  x"4c",  x"2c",  x"4f",  x"2c",  x"50", -- 0420
         x"2c",  x"53",  x"29",  x"3f",  x"20",  x"3a",  x"00",  x"01", -- 0428
         x"27",  x"19",  x"cd",  x"7a",  x"c5",  x"eb",  x"06",  x"0f", -- 0430
         x"1a",  x"13",  x"c5",  x"01",  x"08",  x"00",  x"21",  x"66", -- 0438
         x"c4",  x"ed",  x"b1",  x"21",  x"6d",  x"00",  x"20",  x"09", -- 0440
         x"0c",  x"3e",  x"80",  x"07",  x"0d",  x"20",  x"fc",  x"b6", -- 0448
         x"77",  x"c1",  x"10",  x"e4",  x"cd",  x"03",  x"f0",  x"2c", -- 0450
         x"cd",  x"03",  x"f0",  x"2c",  x"2a",  x"46",  x"00",  x"2b", -- 0458
         x"36",  x"0d",  x"23",  x"c3",  x"f8",  x"c8",  x"32",  x"4f", -- 0460
         x"42",  x"ff",  x"53",  x"2b",  x"50",  x"4c",  x"dd",  x"dd", -- 0468
         x"46",  x"49",  x"4e",  x"44",  x"01",  x"cd",  x"03",  x"f0", -- 0470
         x"23",  x"54",  x"45",  x"58",  x"54",  x"20",  x"3a",  x"00", -- 0478
         x"01",  x"27",  x"06",  x"cd",  x"7a",  x"c5",  x"da",  x"97", -- 0480
         x"c2",  x"11",  x"4b",  x"00",  x"01",  x"22",  x"00",  x"ed", -- 0488
         x"b0",  x"cd",  x"97",  x"c4",  x"c3",  x"26",  x"c5",  x"3a", -- 0490
         x"49",  x"00",  x"b7",  x"28",  x"06",  x"16",  x"00",  x"5f", -- 0498
         x"cd",  x"87",  x"c7",  x"cd",  x"27",  x"c2",  x"ed",  x"5b", -- 04A0
         x"46",  x"00",  x"2a",  x"42",  x"00",  x"af",  x"ed",  x"52", -- 04A8
         x"28",  x"5a",  x"44",  x"4d",  x"eb",  x"11",  x"4b",  x"00", -- 04B0
         x"1a",  x"b7",  x"c8",  x"ed",  x"b1",  x"20",  x"4d",  x"e5", -- 04B8
         x"c5",  x"13",  x"1a",  x"b7",  x"28",  x"08",  x"ed",  x"a1", -- 04C0
         x"28",  x"f7",  x"c1",  x"e1",  x"18",  x"e7",  x"c1",  x"d1", -- 04C8
         x"ed",  x"5b",  x"46",  x"00",  x"2b",  x"ed",  x"52",  x"c8", -- 04D0
         x"44",  x"4d",  x"ed",  x"5b",  x"44",  x"00",  x"2a",  x"46", -- 04D8
         x"00",  x"ed",  x"b0",  x"ed",  x"53",  x"44",  x"00",  x"22", -- 04E0
         x"46",  x"00",  x"11",  x"01",  x"00",  x"cd",  x"c2",  x"c7", -- 04E8
         x"c9",  x"dd",  x"dd",  x"54",  x"4f",  x"50",  x"01",  x"cd", -- 04F0
         x"27",  x"c2",  x"cd",  x"c2",  x"c7",  x"18",  x"27",  x"dd", -- 04F8
         x"dd",  x"42",  x"4f",  x"54",  x"4f",  x"4d",  x"01",  x"cd", -- 0500
         x"0c",  x"c5",  x"18",  x"1a",  x"11",  x"00",  x"00",  x"cd", -- 0508
         x"87",  x"c7",  x"21",  x"27",  x"1d",  x"22",  x"48",  x"00", -- 0510
         x"11",  x"1b",  x"00",  x"cd",  x"c2",  x"c7",  x"c9",  x"dd", -- 0518
         x"dd",  x"45",  x"44",  x"49",  x"54",  x"01",  x"cd",  x"9f", -- 0520
         x"c1",  x"3e",  x"1f",  x"32",  x"9f",  x"b7",  x"cd",  x"a1", -- 0528
         x"c8",  x"cd",  x"63",  x"c7",  x"fe",  x"03",  x"20",  x"0a", -- 0530
         x"cd",  x"09",  x"c8",  x"20",  x"14",  x"21",  x"de",  x"c0", -- 0538
         x"e3",  x"c9",  x"cd",  x"09",  x"c6",  x"2a",  x"a0",  x"b7", -- 0540
         x"22",  x"48",  x"00",  x"3a",  x"4a",  x"00",  x"b7",  x"28", -- 0548
         x"e0",  x"cd",  x"55",  x"c7",  x"18",  x"d8",  x"cd",  x"03", -- 0550
         x"f0",  x"23",  x"20",  x"28",  x"59",  x"2f",  x"4e",  x"20", -- 0558
         x"3f",  x"29",  x"00",  x"cd",  x"63",  x"c7",  x"fe",  x"59", -- 0560
         x"28",  x"05",  x"fe",  x"4e",  x"20",  x"f5",  x"37",  x"f5", -- 0568
         x"cd",  x"03",  x"f0",  x"24",  x"cd",  x"03",  x"f0",  x"2c", -- 0570
         x"f1",  x"c9",  x"cd",  x"63",  x"c7",  x"ed",  x"5b",  x"a0", -- 0578
         x"b7",  x"cd",  x"03",  x"f0",  x"32",  x"fe",  x"03",  x"37", -- 0580
         x"c8",  x"fe",  x"02",  x"28",  x"ed",  x"fe",  x"0c",  x"28", -- 0588
         x"e9",  x"fe",  x"1a",  x"28",  x"e5",  x"fe",  x"11",  x"28", -- 0590
         x"e1",  x"fe",  x"12",  x"28",  x"dd",  x"fe",  x"0a",  x"28", -- 0598
         x"d9",  x"fe",  x"0d",  x"28",  x"1f",  x"fe",  x"05",  x"20", -- 05A0
         x"03",  x"3e",  x"09",  x"77",  x"cd",  x"03",  x"f0",  x"24", -- 05A8
         x"3a",  x"a0",  x"b7",  x"b8",  x"38",  x"06",  x"b9",  x"38", -- 05B0
         x"04",  x"79",  x"18",  x"01",  x"78",  x"5f",  x"ed",  x"53", -- 05B8
         x"a0",  x"b7",  x"18",  x"b6",  x"58",  x"cd",  x"03",  x"f0", -- 05C0
         x"32",  x"a7",  x"c9",  x"cd",  x"03",  x"f0",  x"23",  x"4e", -- 05C8
         x"41",  x"4d",  x"45",  x"20",  x"3a",  x"00",  x"01",  x"0d", -- 05D0
         x"06",  x"78",  x"32",  x"a0",  x"b7",  x"cd",  x"7a",  x"c5", -- 05D8
         x"3e",  x"0e",  x"32",  x"a0",  x"b7",  x"c9",  x"cd",  x"cb", -- 05E0
         x"c5",  x"d8",  x"cd",  x"03",  x"f0",  x"23",  x"41",  x"53", -- 05E8
         x"4d",  x"0d",  x"0a",  x"00",  x"3a",  x"a1",  x"b7",  x"3d", -- 05F0
         x"57",  x"cd",  x"03",  x"f0",  x"32",  x"c9",  x"21",  x"00", -- 05F8
         x"b7",  x"06",  x"80",  x"36",  x"00",  x"23",  x"10",  x"fb", -- 0600
         x"c9",  x"fe",  x"01",  x"ca",  x"c7",  x"c6",  x"fe",  x"08", -- 0608
         x"ca",  x"c7",  x"c6",  x"fe",  x"09",  x"ca",  x"e9",  x"c6", -- 0610
         x"fe",  x"05",  x"ca",  x"a8",  x"c6",  x"fe",  x"0b",  x"28", -- 0618
         x"65",  x"fe",  x"0a",  x"28",  x"48",  x"fe",  x"0d",  x"ca", -- 0620
         x"05",  x"c7",  x"fe",  x"11",  x"28",  x"32",  x"fe",  x"12", -- 0628
         x"28",  x"15",  x"fe",  x"06",  x"ca",  x"41",  x"c7",  x"fe", -- 0630
         x"20",  x"30",  x"51",  x"21",  x"9f",  x"b7",  x"36",  x"1e", -- 0638
         x"cd",  x"03",  x"f0",  x"24",  x"36",  x"1f",  x"c9",  x"cd", -- 0640
         x"09",  x"c8",  x"c0",  x"11",  x"1a",  x"00",  x"cd",  x"87", -- 0648
         x"c7",  x"2a",  x"42",  x"00",  x"ed",  x"5b",  x"46",  x"00", -- 0650
         x"ed",  x"52",  x"cc",  x"12",  x"c5",  x"c3",  x"a1",  x"c8", -- 0658
         x"cd",  x"09",  x"c8",  x"c0",  x"11",  x"1b",  x"00",  x"cd", -- 0660
         x"c2",  x"c7",  x"c3",  x"a1",  x"c8",  x"cd",  x"86",  x"c6", -- 0668
         x"7c",  x"fe",  x"1e",  x"c0",  x"2a",  x"46",  x"00",  x"7e", -- 0670
         x"fe",  x"03",  x"c8",  x"cd",  x"22",  x"c7",  x"3a",  x"4a", -- 0678
         x"00",  x"b7",  x"c0",  x"c3",  x"c0",  x"c8",  x"cd",  x"03", -- 0680
         x"f0",  x"24",  x"3e",  x"0d",  x"2a",  x"a0",  x"b7",  x"cd", -- 0688
         x"03",  x"f0",  x"24",  x"3a",  x"a1",  x"b7",  x"bc",  x"28", -- 0690
         x"06",  x"2e",  x"27",  x"22",  x"a0",  x"b7",  x"c9",  x"fe", -- 0698
         x"1e",  x"20",  x"01",  x"3d",  x"32",  x"a1",  x"b7",  x"c9", -- 06A0
         x"3a",  x"a0",  x"b7",  x"2f",  x"e6",  x"07",  x"3c",  x"47", -- 06A8
         x"d5",  x"3e",  x"1a",  x"cd",  x"8c",  x"c6",  x"54",  x"5d", -- 06B0
         x"cd",  x"03",  x"f0",  x"32",  x"36",  x"00",  x"3e",  x"09", -- 06B8
         x"cd",  x"8c",  x"c6",  x"10",  x"ec",  x"d1",  x"c9",  x"47", -- 06C0
         x"cd",  x"03",  x"f0",  x"24",  x"ed",  x"5b",  x"a0",  x"b7", -- 06C8
         x"7b",  x"fe",  x"27",  x"20",  x"04",  x"3e",  x"09",  x"18", -- 06D0
         x"ef",  x"e6",  x"07",  x"c8",  x"cd",  x"03",  x"f0",  x"32", -- 06D8
         x"af",  x"be",  x"c0",  x"2b",  x"be",  x"78",  x"28",  x"e0", -- 06E0
         x"c9",  x"3e",  x"09",  x"cd",  x"8c",  x"c6",  x"ed",  x"5b", -- 06E8
         x"a0",  x"b7",  x"7b",  x"fe",  x"27",  x"c8",  x"e6",  x"07", -- 06F0
         x"c8",  x"cd",  x"03",  x"f0",  x"32",  x"af",  x"be",  x"c0", -- 06F8
         x"2b",  x"be",  x"28",  x"e5",  x"c9",  x"3a",  x"a1",  x"b7", -- 0700
         x"fe",  x"1d",  x"28",  x"16",  x"3c",  x"57",  x"1e",  x"00", -- 0708
         x"cd",  x"03",  x"f0",  x"32",  x"06",  x"28",  x"af",  x"be", -- 0710
         x"20",  x"08",  x"23",  x"10",  x"fa",  x"3e",  x"0a",  x"c3", -- 0718
         x"6d",  x"c6",  x"21",  x"28",  x"b2",  x"cd",  x"2a",  x"c8", -- 0720
         x"3a",  x"a1",  x"b7",  x"3c",  x"32",  x"9f",  x"b7",  x"3e", -- 0728
         x"0d",  x"cd",  x"03",  x"f0",  x"24",  x"3e",  x"0a",  x"cd", -- 0730
         x"03",  x"f0",  x"24",  x"3e",  x"1f",  x"32",  x"9f",  x"b7", -- 0738
         x"c9",  x"3a",  x"4b",  x"00",  x"b7",  x"c8",  x"cd",  x"09", -- 0740
         x"c8",  x"11",  x"01",  x"00",  x"cd",  x"87",  x"c7",  x"cd", -- 0748
         x"97",  x"c4",  x"c3",  x"a1",  x"c8",  x"2a",  x"a0",  x"b7", -- 0750
         x"3e",  x"1d",  x"32",  x"a1",  x"b7",  x"cd",  x"6a",  x"c7", -- 0758
         x"22",  x"a0",  x"b7",  x"c5",  x"cd",  x"03",  x"f0",  x"04", -- 0760
         x"c1",  x"c9",  x"cd",  x"03",  x"f0",  x"23",  x"0d",  x"3e", -- 0768
         x"3e",  x"3e",  x"20",  x"4e",  x"4f",  x"20",  x"4d",  x"45", -- 0770
         x"4d",  x"4f",  x"52",  x"59",  x"20",  x"3c",  x"3c",  x"3c", -- 0778
         x"0a",  x"00",  x"af",  x"32",  x"4a",  x"00",  x"c9",  x"2a", -- 0780
         x"42",  x"00",  x"ed",  x"4b",  x"46",  x"00",  x"c5",  x"af", -- 0788
         x"ed",  x"42",  x"44",  x"4d",  x"e1",  x"c8",  x"3e",  x"0d", -- 0790
         x"ed",  x"b1",  x"e2",  x"a8",  x"c7",  x"1b",  x"7a",  x"b3", -- 0798
         x"20",  x"f4",  x"7e",  x"fe",  x"0a",  x"20",  x"01",  x"23", -- 07A0
         x"ed",  x"5b",  x"46",  x"00",  x"d5",  x"af",  x"ed",  x"52", -- 07A8
         x"44",  x"4d",  x"e1",  x"c8",  x"ed",  x"5b",  x"44",  x"00", -- 07B0
         x"ed",  x"b0",  x"ed",  x"53",  x"44",  x"00",  x"22",  x"46", -- 07B8
         x"00",  x"c9",  x"2a",  x"44",  x"00",  x"ed",  x"4b",  x"40", -- 07C0
         x"00",  x"e5",  x"af",  x"ed",  x"42",  x"44",  x"4d",  x"e1", -- 07C8
         x"c8",  x"2b",  x"3e",  x"0d",  x"ed",  x"b9",  x"e2",  x"df", -- 07D0
         x"c7",  x"1b",  x"7a",  x"b3",  x"20",  x"f4",  x"23",  x"23", -- 07D8
         x"7e",  x"fe",  x"0a",  x"20",  x"01",  x"23",  x"eb",  x"2a", -- 07E0
         x"44",  x"00",  x"e5",  x"af",  x"ed",  x"52",  x"44",  x"4d", -- 07E8
         x"e1",  x"28",  x"11",  x"ed",  x"5b",  x"46",  x"00",  x"1b", -- 07F0
         x"2b",  x"ed",  x"b8",  x"13",  x"ed",  x"53",  x"46",  x"00", -- 07F8
         x"23",  x"22",  x"44",  x"00",  x"3a",  x"4a",  x"00",  x"b7", -- 0800
         x"c9",  x"2a",  x"44",  x"00",  x"e5",  x"21",  x"28",  x"b2", -- 0808
         x"11",  x"28",  x"00",  x"06",  x"1e",  x"c5",  x"d5",  x"e5", -- 0810
         x"cd",  x"2a",  x"c8",  x"e1",  x"d1",  x"c1",  x"3a",  x"4a", -- 0818
         x"00",  x"b7",  x"20",  x"03",  x"19",  x"10",  x"ee",  x"d1", -- 0820
         x"18",  x"bd",  x"54",  x"5d",  x"01",  x"28",  x"00",  x"09", -- 0828
         x"2b",  x"03",  x"af",  x"ed",  x"a9",  x"e0",  x"28",  x"fb", -- 0830
         x"d5",  x"e5",  x"2a",  x"46",  x"00",  x"ed",  x"5b",  x"44", -- 0838
         x"00",  x"2b",  x"2b",  x"37",  x"ed",  x"52",  x"e1",  x"d1", -- 0840
         x"30",  x"06",  x"3e",  x"01",  x"32",  x"4a",  x"00",  x"c9", -- 0848
         x"03",  x"23",  x"7e",  x"fe",  x"21",  x"30",  x"10",  x"ed", -- 0850
         x"a9",  x"e2",  x"60",  x"c8",  x"28",  x"f9",  x"18",  x"f0", -- 0858
         x"06",  x"01",  x"3e",  x"20",  x"12",  x"18",  x"04",  x"23", -- 0860
         x"ed",  x"52",  x"45",  x"2a",  x"44",  x"00",  x"eb",  x"7e", -- 0868
         x"b7",  x"20",  x"0e",  x"0e",  x"08",  x"23",  x"05",  x"0d", -- 0870
         x"28",  x"03",  x"be",  x"28",  x"f8",  x"04",  x"2b",  x"3e", -- 0878
         x"09",  x"e5",  x"2a",  x"46",  x"00",  x"2b",  x"37",  x"ed", -- 0880
         x"52",  x"e1",  x"20",  x"05",  x"cd",  x"4a",  x"c8",  x"18", -- 0888
         x"05",  x"12",  x"13",  x"23",  x"10",  x"d9",  x"eb",  x"36", -- 0890
         x"0d",  x"23",  x"36",  x"0a",  x"23",  x"22",  x"44",  x"00", -- 0898
         x"c9",  x"cd",  x"03",  x"f0",  x"2d",  x"0e",  x"1e",  x"3e", -- 08A0
         x"02",  x"cd",  x"03",  x"f0",  x"24",  x"cd",  x"c0",  x"c8", -- 08A8
         x"3e",  x"0a",  x"cd",  x"03",  x"f0",  x"24",  x"0d",  x"20", -- 08B0
         x"ee",  x"2a",  x"48",  x"00",  x"22",  x"a0",  x"b7",  x"c9", -- 08B8
         x"ed",  x"5b",  x"46",  x"00",  x"1a",  x"fe",  x"03",  x"c8", -- 08C0
         x"fe",  x"09",  x"20",  x"05",  x"cd",  x"a8",  x"c6",  x"18", -- 08C8
         x"03",  x"cd",  x"8c",  x"c6",  x"1a",  x"13",  x"fe",  x"0d", -- 08D0
         x"20",  x"ea",  x"1a",  x"fe",  x"0a",  x"20",  x"01",  x"13", -- 08D8
         x"ed",  x"53",  x"46",  x"00",  x"1a",  x"fe",  x"03",  x"c0", -- 08E0
         x"2a",  x"48",  x"00",  x"ed",  x"5b",  x"a0",  x"b7",  x"14", -- 08E8
         x"ed",  x"52",  x"d8",  x"ed",  x"53",  x"48",  x"00",  x"c9", -- 08F0
         x"e5",  x"21",  x"6d",  x"00",  x"cb",  x"56",  x"20",  x"06", -- 08F8
         x"2a",  x"72",  x"00",  x"22",  x"74",  x"00",  x"c3",  x"6d", -- 0900
         x"ca",  x"7e",  x"fe",  x"20",  x"28",  x"03",  x"fe",  x"09", -- 0908
         x"c0",  x"23",  x"18",  x"f5",  x"7e",  x"fe",  x"20",  x"30", -- 0910
         x"25",  x"23",  x"e5",  x"d5",  x"c5",  x"23",  x"13",  x"1a", -- 0918
         x"cd",  x"40",  x"c9",  x"38",  x"0a",  x"47",  x"7e",  x"cd", -- 0920
         x"40",  x"c9",  x"b8",  x"20",  x"0d",  x"18",  x"ee",  x"7e", -- 0928
         x"cd",  x"40",  x"c9",  x"30",  x"05",  x"c1",  x"e1",  x"e1", -- 0930
         x"b7",  x"c9",  x"c1",  x"d1",  x"e1",  x"2b",  x"37",  x"c9", -- 0938
         x"cd",  x"de",  x"d1",  x"d0",  x"fe",  x"30",  x"38",  x"04", -- 0940
         x"fe",  x"3a",  x"3f",  x"d0",  x"fe",  x"2e",  x"c8",  x"fe", -- 0948
         x"5f",  x"c8",  x"37",  x"c9",  x"3a",  x"88",  x"00",  x"fe", -- 0950
         x"20",  x"28",  x"16",  x"3e",  x"2a",  x"32",  x"89",  x"00", -- 0958
         x"2a",  x"7c",  x"00",  x"7d",  x"3c",  x"27",  x"6f",  x"30", -- 0960
         x"05",  x"af",  x"7c",  x"3c",  x"27",  x"67",  x"22",  x"7c", -- 0968
         x"00",  x"21",  x"88",  x"00",  x"11",  x"40",  x"00",  x"3a", -- 0970
         x"6d",  x"00",  x"e6",  x"20",  x"28",  x"02",  x"1e",  x"27", -- 0978
         x"7e",  x"23",  x"fe",  x"0d",  x"28",  x"07",  x"cd",  x"ef", -- 0980
         x"d1",  x"7b",  x"b7",  x"20",  x"f3",  x"3e",  x"0d",  x"cd", -- 0988
         x"ef",  x"d1",  x"3e",  x"0a",  x"cd",  x"ef",  x"d1",  x"21", -- 0990
         x"88",  x"00",  x"54",  x"5d",  x"13",  x"01",  x"40",  x"00", -- 0998
         x"36",  x"20",  x"ed",  x"b0",  x"36",  x"0d",  x"c9",  x"21", -- 09A0
         x"8a",  x"00",  x"7a",  x"cd",  x"af",  x"c9",  x"7b",  x"f5", -- 09A8
         x"1f",  x"1f",  x"1f",  x"1f",  x"cd",  x"b8",  x"c9",  x"f1", -- 09B0
         x"e6",  x"0f",  x"c6",  x"30",  x"fe",  x"3a",  x"38",  x"02", -- 09B8
         x"c6",  x"07",  x"77",  x"23",  x"c9",  x"cd",  x"93",  x"ca", -- 09C0
         x"3a",  x"6d",  x"00",  x"17",  x"30",  x"3e",  x"e5",  x"f5", -- 09C8
         x"1f",  x"1f",  x"dc",  x"54",  x"c9",  x"f1",  x"cb",  x"6f", -- 09D0
         x"f5",  x"20",  x"08",  x"3a",  x"88",  x"00",  x"fe",  x"20", -- 09D8
         x"c4",  x"54",  x"c9",  x"cd",  x"97",  x"c9",  x"cd",  x"03", -- 09E0
         x"f0",  x"2a",  x"30",  x"06",  x"f1",  x"e1",  x"20",  x"5a", -- 09E8
         x"e1",  x"c9",  x"f1",  x"ed",  x"5b",  x"7a",  x"00",  x"cd", -- 09F0
         x"a7",  x"c9",  x"23",  x"22",  x"76",  x"00",  x"e1",  x"e5", -- 09F8
         x"11",  x"98",  x"00",  x"01",  x"30",  x"00",  x"ed",  x"b0", -- 0A00
         x"eb",  x"36",  x"0d",  x"e1",  x"7e",  x"fe",  x"03",  x"20", -- 0A08
         x"b4",  x"cd",  x"97",  x"c9",  x"21",  x"6d",  x"00",  x"7e", -- 0A10
         x"17",  x"30",  x"3c",  x"e6",  x"20",  x"20",  x"2b",  x"cd", -- 0A18
         x"03",  x"f0",  x"23",  x"0a",  x"45",  x"52",  x"52",  x"4f", -- 0A20
         x"52",  x"53",  x"3a",  x"20",  x"00",  x"2a",  x"7c",  x"00", -- 0A28
         x"cd",  x"03",  x"f0",  x"1a",  x"cd",  x"03",  x"f0",  x"23", -- 0A30
         x"0d",  x"0a",  x"0a",  x"00",  x"21",  x"6d",  x"00",  x"cb", -- 0A38
         x"5e",  x"28",  x"12",  x"36",  x"98",  x"cd",  x"2e",  x"d2", -- 0A40
         x"18",  x"21",  x"01",  x"a0",  x"00",  x"cd",  x"03",  x"f0", -- 0A48
         x"09",  x"cd",  x"03",  x"f0",  x"2c",  x"e1",  x"c9",  x"cb", -- 0A50
         x"fe",  x"cd",  x"03",  x"f0",  x"23",  x"45",  x"4e",  x"44", -- 0A58
         x"20",  x"50",  x"41",  x"53",  x"53",  x"20",  x"31",  x"0d", -- 0A60
         x"0a",  x"0a",  x"00",  x"e1",  x"e5",  x"21",  x"00",  x"00", -- 0A68
         x"22",  x"7c",  x"00",  x"22",  x"7e",  x"00",  x"3a",  x"6d", -- 0A70
         x"00",  x"e6",  x"82",  x"fe",  x"82",  x"20",  x"07",  x"21", -- 0A78
         x"00",  x"c4",  x"cd",  x"03",  x"f0",  x"1e",  x"e1",  x"e5", -- 0A80
         x"fd",  x"2a",  x"70",  x"00",  x"fd",  x"22",  x"7a",  x"00", -- 0A88
         x"c3",  x"c8",  x"c9",  x"0e",  x"ff",  x"cd",  x"de",  x"d1", -- 0A90
         x"30",  x"18",  x"cd",  x"09",  x"c9",  x"fe",  x"0d",  x"28", -- 0A98
         x"0e",  x"fe",  x"3b",  x"28",  x"0a",  x"cd",  x"de",  x"d1", -- 0AA0
         x"30",  x"48",  x"3e",  x"31",  x"32",  x"88",  x"00",  x"c3", -- 0AA8
         x"a6",  x"cb",  x"0c",  x"54",  x"5d",  x"cd",  x"1a",  x"c9", -- 0AB0
         x"eb",  x"fe",  x"3a",  x"20",  x"01",  x"23",  x"3a",  x"6d", -- 0AB8
         x"00",  x"17",  x"38",  x"d6",  x"eb",  x"d5",  x"cd",  x"1a", -- 0AC0
         x"d0",  x"d1",  x"38",  x"06",  x"2b",  x"36",  x"01",  x"eb", -- 0AC8
         x"18",  x"c8",  x"d5",  x"eb",  x"3e",  x"3a",  x"2b",  x"be", -- 0AD0
         x"20",  x"05",  x"7e",  x"cd",  x"de",  x"d1",  x"2b",  x"12", -- 0AD8
         x"1b",  x"fe",  x"20",  x"30",  x"f5",  x"2a",  x"7a",  x"00", -- 0AE0
         x"eb",  x"72",  x"2b",  x"73",  x"22",  x"74",  x"00",  x"e1", -- 0AE8
         x"18",  x"a8",  x"11",  x"00",  x"00",  x"d6",  x"40",  x"47", -- 0AF0
         x"83",  x"5f",  x"7a",  x"82",  x"80",  x"57",  x"23",  x"7e", -- 0AF8
         x"cd",  x"de",  x"d1",  x"30",  x"f0",  x"e5",  x"fe",  x"20", -- 0B00
         x"28",  x"0c",  x"fe",  x"09",  x"28",  x"08",  x"fe",  x"3b", -- 0B08
         x"28",  x"04",  x"fe",  x"0d",  x"20",  x"5a",  x"a7",  x"21", -- 0B10
         x"2b",  x"4b",  x"ed",  x"52",  x"28",  x"18",  x"7a",  x"01", -- 0B18
         x"1d",  x"00",  x"21",  x"a8",  x"d1",  x"ed",  x"b1",  x"20", -- 0B20
         x"2d",  x"3e",  x"03",  x"b9",  x"38",  x"22",  x"7a",  x"83", -- 0B28
         x"fe",  x"73",  x"38",  x"fb",  x"18",  x"e9",  x"79",  x"b7", -- 0B30
         x"3e",  x"37",  x"20",  x"36",  x"e1",  x"cd",  x"3b",  x"cf", -- 0B38
         x"3a",  x"6d",  x"00",  x"17",  x"38",  x"60",  x"e5",  x"2a", -- 0B40
         x"74",  x"00",  x"73",  x"23",  x"72",  x"e1",  x"18",  x"56", -- 0B48
         x"01",  x"1c",  x"00",  x"09",  x"53",  x"5e",  x"7a",  x"16", -- 0B50
         x"00",  x"21",  x"09",  x"d1",  x"19",  x"46",  x"21",  x"50", -- 0B58
         x"d1",  x"19",  x"4e",  x"e6",  x"07",  x"57",  x"79",  x"0f", -- 0B60
         x"0f",  x"0f",  x"0f",  x"e6",  x"07",  x"92",  x"28",  x"05", -- 0B68
         x"3e",  x"34",  x"32",  x"88",  x"00",  x"e1",  x"20",  x"2e", -- 0B70
         x"c5",  x"af",  x"32",  x"78",  x"00",  x"79",  x"fe",  x"4e", -- 0B78
         x"28",  x"17",  x"e5",  x"cd",  x"d8",  x"ce",  x"dc",  x"70", -- 0B80
         x"ce",  x"2b",  x"7e",  x"23",  x"fe",  x"2c",  x"cc",  x"70", -- 0B88
         x"ce",  x"3a",  x"78",  x"00",  x"b7",  x"c4",  x"9f",  x"ce", -- 0B90
         x"e1",  x"f1",  x"f5",  x"3e",  x"ed",  x"fc",  x"9f",  x"ce", -- 0B98
         x"3e",  x"0f",  x"c1",  x"cd",  x"ba",  x"cb",  x"fd",  x"22", -- 0BA0
         x"7a",  x"00",  x"3e",  x"0d",  x"c5",  x"01",  x"00",  x"01", -- 0BA8
         x"ed",  x"b1",  x"7e",  x"fe",  x"0a",  x"20",  x"01",  x"23", -- 0BB0
         x"c1",  x"c9",  x"e5",  x"c5",  x"a1",  x"21",  x"d2",  x"cb", -- 0BB8
         x"11",  x"2b",  x"cf",  x"3c",  x"06",  x"00",  x"f5",  x"1a", -- 0BC0
         x"13",  x"4f",  x"09",  x"f1",  x"3d",  x"20",  x"f7",  x"c1", -- 0BC8
         x"e3",  x"c9",  x"3e",  x"cb",  x"cd",  x"9f",  x"ce",  x"3a", -- 0BD0
         x"82",  x"00",  x"b7",  x"28",  x"06",  x"3a",  x"80",  x"00", -- 0BD8
         x"cd",  x"9f",  x"ce",  x"cd",  x"70",  x"ce",  x"7b",  x"07", -- 0BE0
         x"07",  x"07",  x"80",  x"f5",  x"cd",  x"70",  x"ce",  x"20", -- 0BE8
         x"02",  x"7b",  x"3d",  x"c1",  x"c3",  x"9b",  x"ce",  x"e5", -- 0BF0
         x"af",  x"32",  x"78",  x"00",  x"cd",  x"70",  x"ce",  x"28", -- 0BF8
         x"20",  x"4f",  x"cd",  x"70",  x"ce",  x"28",  x"50",  x"5f", -- 0C00
         x"81",  x"fe",  x"0f",  x"d2",  x"c6",  x"cc",  x"e1",  x"7b", -- 0C08
         x"c6",  x"40",  x"47",  x"79",  x"cd",  x"98",  x"ce",  x"3a", -- 0C10
         x"78",  x"00",  x"b7",  x"c8",  x"3a",  x"79",  x"00",  x"18", -- 0C18
         x"47",  x"d1",  x"3a",  x"87",  x"00",  x"3c",  x"28",  x"03", -- 0C20
         x"3c",  x"18",  x"3d",  x"ed",  x"4b",  x"80",  x"00",  x"cd", -- 0C28
         x"70",  x"ce",  x"ed",  x"43",  x"80",  x"00",  x"fe",  x"07", -- 0C30
         x"20",  x"07",  x"3e",  x"32",  x"cd",  x"9f",  x"ce",  x"18", -- 0C38
         x"44",  x"fe",  x"20",  x"06",  x"22",  x"28",  x"0a",  x"f5", -- 0C40
         x"3e",  x"ed",  x"cd",  x"9f",  x"ce",  x"f1",  x"c6",  x"43", -- 0C48
         x"47",  x"78",  x"cd",  x"9f",  x"ce",  x"18",  x"2e",  x"e1", -- 0C50
         x"fe",  x"28",  x"20",  x"10",  x"32",  x"78",  x"00",  x"3a", -- 0C58
         x"87",  x"00",  x"fe",  x"ff",  x"28",  x"06",  x"c6",  x"0a", -- 0C60
         x"cd",  x"9f",  x"ce",  x"c9",  x"cd",  x"3b",  x"cf",  x"3a", -- 0C68
         x"87",  x"00",  x"fe",  x"07",  x"20",  x"12",  x"3a",  x"78", -- 0C70
         x"00",  x"fe",  x"28",  x"20",  x"0b",  x"3e",  x"3a",  x"cd", -- 0C78
         x"9f",  x"ce",  x"cd",  x"3b",  x"cf",  x"c3",  x"8e",  x"ce", -- 0C80
         x"fe",  x"06",  x"28",  x"0a",  x"3a",  x"86",  x"00",  x"fe", -- 0C88
         x"12",  x"3a",  x"87",  x"00",  x"30",  x"0e",  x"06",  x"06", -- 0C90
         x"cd",  x"98",  x"ce",  x"cd",  x"18",  x"cd",  x"cd",  x"3b", -- 0C98
         x"cf",  x"7b",  x"18",  x"c4",  x"f5",  x"cd",  x"70",  x"ce", -- 0CA0
         x"fe",  x"28",  x"0e",  x"01",  x"20",  x"11",  x"0e",  x"4b", -- 0CA8
         x"f1",  x"f5",  x"fe",  x"20",  x"20",  x"04",  x"0e",  x"0a", -- 0CB0
         x"18",  x"05",  x"3e",  x"ed",  x"cd",  x"9f",  x"ce",  x"79", -- 0CB8
         x"c1",  x"cd",  x"9b",  x"ce",  x"18",  x"bf",  x"e1",  x"cd", -- 0CC0
         x"70",  x"ce",  x"fe",  x"30",  x"20",  x"04",  x"3e",  x"f9", -- 0CC8
         x"18",  x"d0",  x"fe",  x"07",  x"20",  x"05",  x"cd",  x"70", -- 0CD0
         x"ce",  x"c6",  x"10",  x"f5",  x"3e",  x"ed",  x"cd",  x"9f", -- 0CD8
         x"ce",  x"f1",  x"18",  x"be",  x"c5",  x"c3",  x"ec",  x"cb", -- 0CE0
         x"cd",  x"70",  x"ce",  x"20",  x"09",  x"3e",  x"46",  x"80", -- 0CE8
         x"cd",  x"9f",  x"ce",  x"7b",  x"18",  x"ec",  x"fe",  x"06", -- 0CF0
         x"28",  x"07",  x"3a",  x"86",  x"00",  x"fe",  x"0c",  x"30", -- 0CF8
         x"21",  x"2b",  x"7e",  x"23",  x"fe",  x"2c",  x"28",  x"e0", -- 0D00
         x"3e",  x"05",  x"b8",  x"3a",  x"87",  x"00",  x"38",  x"05", -- 0D08
         x"cd",  x"98",  x"ce",  x"18",  x"03",  x"cd",  x"9b",  x"ce", -- 0D10
         x"3a",  x"82",  x"00",  x"b7",  x"c8",  x"3a",  x"80",  x"00", -- 0D18
         x"18",  x"c0",  x"eb",  x"21",  x"43",  x"cd",  x"78",  x"ed", -- 0D20
         x"b1",  x"46",  x"eb",  x"2b",  x"7e",  x"23",  x"fe",  x"2c", -- 0D28
         x"3a",  x"87",  x"00",  x"c2",  x"9b",  x"ce",  x"78",  x"fe", -- 0D30
         x"40",  x"38",  x"a9",  x"c5",  x"3e",  x"ed",  x"cd",  x"9f", -- 0D38
         x"ce",  x"18",  x"a2",  x"05",  x"0b",  x"04",  x"03",  x"80", -- 0D40
         x"09",  x"88",  x"4a",  x"98",  x"42",  x"cd",  x"3b",  x"cf", -- 0D48
         x"7b",  x"11",  x"59",  x"cd",  x"83",  x"5f",  x"1a",  x"18", -- 0D50
         x"17",  x"46",  x"56",  x"5e",  x"cd",  x"70",  x"ce",  x"4f", -- 0D58
         x"cd",  x"70",  x"ce",  x"3a",  x"87",  x"00",  x"fe",  x"ff", -- 0D60
         x"20",  x"0b",  x"3e",  x"db",  x"cd",  x"9f",  x"ce",  x"7b", -- 0D68
         x"cd",  x"9f",  x"ce",  x"c9",  x"4b",  x"3e",  x"ed",  x"cd", -- 0D70
         x"9f",  x"ce",  x"79",  x"c3",  x"98",  x"ce",  x"cd",  x"70", -- 0D78
         x"ce",  x"3a",  x"87",  x"00",  x"fe",  x"ff",  x"f5",  x"4b", -- 0D80
         x"cd",  x"70",  x"ce",  x"5f",  x"f1",  x"20",  x"e5",  x"3e", -- 0D88
         x"d3",  x"cd",  x"9f",  x"ce",  x"79",  x"18",  x"89",  x"3e", -- 0D90
         x"cb",  x"cd",  x"9f",  x"ce",  x"cd",  x"70",  x"ce",  x"80", -- 0D98
         x"47",  x"3a",  x"82",  x"00",  x"b7",  x"28",  x"04",  x"7b", -- 0DA0
         x"cd",  x"9f",  x"ce",  x"18",  x"1a",  x"cd",  x"70",  x"ce", -- 0DA8
         x"06",  x"e3",  x"fe",  x"28",  x"28",  x"11",  x"06",  x"eb", -- 0DB0
         x"fe",  x"10",  x"28",  x"0b",  x"06",  x"08",  x"fe",  x"30", -- 0DB8
         x"28",  x"05",  x"3e",  x"39",  x"c3",  x"56",  x"ce",  x"c3", -- 0DC0
         x"9e",  x"ce",  x"cd",  x"d8",  x"ce",  x"30",  x"14",  x"cd", -- 0DC8
         x"70",  x"ce",  x"28",  x"18",  x"3a",  x"86",  x"00",  x"fe", -- 0DD0
         x"3a",  x"06",  x"e9",  x"28",  x"ea",  x"3e",  x"41",  x"32", -- 0DD8
         x"88",  x"00",  x"c9",  x"cd",  x"98",  x"ce",  x"cd",  x"3b", -- 0DE0
         x"cf",  x"c3",  x"8e",  x"ce",  x"78",  x"06",  x"c3",  x"fe", -- 0DE8
         x"c2",  x"28",  x"02",  x"06",  x"cd",  x"78",  x"c3",  x"3c", -- 0DF0
         x"cc",  x"cd",  x"d8",  x"ce",  x"d2",  x"98",  x"ce",  x"cd", -- 0DF8
         x"70",  x"ce",  x"3a",  x"84",  x"00",  x"b7",  x"20",  x"d5", -- 0E00
         x"3e",  x"c9",  x"c3",  x"9f",  x"ce",  x"cd",  x"d8",  x"ce", -- 0E08
         x"30",  x"07",  x"cd",  x"70",  x"ce",  x"20",  x"c6",  x"18", -- 0E10
         x"23",  x"06",  x"20",  x"cd",  x"98",  x"ce",  x"cd",  x"3b", -- 0E18
         x"cf",  x"e5",  x"fd",  x"e5",  x"eb",  x"d1",  x"37",  x"ed", -- 0E20
         x"52",  x"5d",  x"7c",  x"cb",  x"03",  x"ce",  x"00",  x"28", -- 0E28
         x"05",  x"3e",  x"36",  x"32",  x"88",  x"00",  x"7d",  x"e1", -- 0E30
         x"cd",  x"9f",  x"ce",  x"c9",  x"78",  x"cd",  x"9f",  x"ce", -- 0E38
         x"18",  x"df",  x"cd",  x"70",  x"ce",  x"7b",  x"cd",  x"9f", -- 0E40
         x"ce",  x"7a",  x"10",  x"fa",  x"c9",  x"cd",  x"09",  x"c9", -- 0E48
         x"fe",  x"27",  x"28",  x"06",  x"3e",  x"38",  x"32",  x"88", -- 0E50
         x"00",  x"c9",  x"23",  x"7e",  x"fe",  x"20",  x"38",  x"f4", -- 0E58
         x"23",  x"fe",  x"27",  x"c8",  x"cd",  x"9f",  x"ce",  x"18", -- 0E60
         x"f2",  x"cd",  x"3b",  x"cf",  x"d5",  x"fd",  x"e1",  x"c9", -- 0E68
         x"cd",  x"3b",  x"cf",  x"3a",  x"82",  x"00",  x"b7",  x"28", -- 0E70
         x"09",  x"32",  x"78",  x"00",  x"3a",  x"80",  x"00",  x"32", -- 0E78
         x"79",  x"00",  x"3a",  x"83",  x"00",  x"fe",  x"28",  x"c8", -- 0E80
         x"3a",  x"87",  x"00",  x"fe",  x"ff",  x"c9",  x"ed",  x"4b", -- 0E88
         x"80",  x"00",  x"79",  x"cd",  x"9f",  x"ce",  x"18",  x"06", -- 0E90
         x"07",  x"07",  x"07",  x"80",  x"18",  x"01",  x"78",  x"d9", -- 0E98
         x"4f",  x"3a",  x"6d",  x"00",  x"17",  x"17",  x"30",  x"08", -- 0EA0
         x"2a",  x"6e",  x"00",  x"fd",  x"e5",  x"d1",  x"19",  x"71", -- 0EA8
         x"1f",  x"30",  x"21",  x"2a",  x"7e",  x"00",  x"23",  x"22", -- 0EB0
         x"7e",  x"00",  x"cb",  x"6f",  x"28",  x"05",  x"cd",  x"54", -- 0EB8
         x"d2",  x"18",  x"11",  x"21",  x"97",  x"00",  x"7d",  x"2a", -- 0EC0
         x"76",  x"00",  x"bd",  x"28",  x"07",  x"79",  x"cd",  x"af", -- 0EC8
         x"c9",  x"22",  x"76",  x"00",  x"d9",  x"fd",  x"23",  x"c9", -- 0ED0
         x"c5",  x"e5",  x"cd",  x"09",  x"c9",  x"cd",  x"de",  x"d1", -- 0ED8
         x"38",  x"35",  x"57",  x"1e",  x"20",  x"23",  x"7e",  x"cd", -- 0EE0
         x"de",  x"d1",  x"38",  x"08",  x"5f",  x"23",  x"7e",  x"cd", -- 0EE8
         x"de",  x"d1",  x"30",  x"23",  x"cd",  x"09",  x"c9",  x"fe", -- 0EF0
         x"2c",  x"20",  x"01",  x"23",  x"e5",  x"21",  x"2a",  x"cf", -- 0EF8
         x"01",  x"10",  x"00",  x"7b",  x"ed",  x"b9",  x"20",  x"0e", -- 0F00
         x"7a",  x"be",  x"20",  x"f7",  x"cb",  x"39",  x"30",  x"06", -- 0F08
         x"79",  x"e1",  x"d1",  x"c1",  x"3f",  x"c9",  x"e1",  x"e1", -- 0F10
         x"c1",  x"37",  x"c9",  x"4e",  x"5a",  x"5a",  x"20",  x"4e", -- 0F18
         x"43",  x"43",  x"20",  x"50",  x"4f",  x"50",  x"45",  x"50", -- 0F20
         x"20",  x"4d",  x"20",  x"00",  x"00",  x"25",  x"ed",  x"04", -- 0F28
         x"65",  x"0f",  x"22",  x"19",  x"16",  x"1d",  x"2f",  x"14", -- 0F30
         x"35",  x"0b",  x"1c",  x"c5",  x"af",  x"d9",  x"06",  x"08", -- 0F38
         x"21",  x"7f",  x"00",  x"23",  x"77",  x"10",  x"fc",  x"35", -- 0F40
         x"d9",  x"3e",  x"2b",  x"32",  x"85",  x"00",  x"18",  x"01", -- 0F48
         x"23",  x"cd",  x"09",  x"c9",  x"7e",  x"fe",  x"3b",  x"28", -- 0F50
         x"30",  x"fe",  x"20",  x"38",  x"2c",  x"32",  x"84",  x"00", -- 0F58
         x"fe",  x"27",  x"ca",  x"f6",  x"cf",  x"fe",  x"2c",  x"28", -- 0F60
         x"1f",  x"fe",  x"28",  x"28",  x"26",  x"fe",  x"29",  x"28", -- 0F68
         x"df",  x"fe",  x"2d",  x"28",  x"23",  x"fe",  x"2b",  x"28", -- 0F70
         x"1f",  x"fe",  x"24",  x"28",  x"04",  x"fe",  x"23",  x"20", -- 0F78
         x"1c",  x"ed",  x"4b",  x"7a",  x"00",  x"c3",  x"16",  x"d0", -- 0F80
         x"23",  x"ed",  x"5b",  x"80",  x"00",  x"c1",  x"3a",  x"84", -- 0F88
         x"00",  x"b7",  x"c9",  x"32",  x"83",  x"00",  x"18",  x"b8", -- 0F90
         x"32",  x"85",  x"00",  x"18",  x"b3",  x"cd",  x"de",  x"d1", -- 0F98
         x"d2",  x"84",  x"d0",  x"e5",  x"0e",  x"0a",  x"cd",  x"d7", -- 0FA0
         x"cf",  x"38",  x"08",  x"e1",  x"23",  x"e5",  x"3e",  x"35", -- 0FA8
         x"32",  x"88",  x"00",  x"0e",  x"10",  x"cd",  x"d7",  x"cf", -- 0FB0
         x"38",  x"fb",  x"e1",  x"fe",  x"11",  x"28",  x"02",  x"0e", -- 0FB8
         x"0a",  x"e5",  x"21",  x"00",  x"00",  x"e3",  x"cd",  x"d7", -- 0FC0
         x"cf",  x"e3",  x"38",  x"1e",  x"fe",  x"11",  x"ca",  x"80", -- 0FC8
         x"d0",  x"e3",  x"2b",  x"e3",  x"c3",  x"80",  x"d0",  x"7e", -- 0FD0
         x"cd",  x"de",  x"d1",  x"23",  x"fe",  x"3a",  x"30",  x"02", -- 0FD8
         x"d6",  x"30",  x"fe",  x"41",  x"38",  x"02",  x"d6",  x"37", -- 0FE0
         x"b9",  x"c9",  x"5f",  x"af",  x"57",  x"19",  x"eb",  x"6f", -- 0FE8
         x"41",  x"19",  x"10",  x"fd",  x"18",  x"cf",  x"01",  x"00", -- 0FF0
         x"00",  x"3a",  x"86",  x"00",  x"fe",  x"2d",  x"ca",  x"50", -- 0FF8
         x"cf",  x"23",  x"7e",  x"fe",  x"27",  x"28",  x"0f",  x"fe", -- 1000
         x"20",  x"38",  x"04",  x"41",  x"4f",  x"18",  x"f2",  x"3e", -- 1008
         x"38",  x"32",  x"88",  x"00",  x"18",  x"01",  x"23",  x"e5", -- 1010
         x"18",  x"44",  x"e5",  x"2a",  x"72",  x"00",  x"e5",  x"ed", -- 1018
         x"5b",  x"74",  x"00",  x"1b",  x"b7",  x"ed",  x"52",  x"44", -- 1020
         x"4d",  x"e1",  x"d1",  x"1a",  x"cd",  x"de",  x"d1",  x"ed", -- 1028
         x"b9",  x"37",  x"e0",  x"cd",  x"14",  x"c9",  x"38",  x"f3", -- 1030
         x"c9",  x"f1",  x"1b",  x"1b",  x"eb",  x"cd",  x"1a",  x"d0", -- 1038
         x"d5",  x"2b",  x"7e",  x"3d",  x"20",  x"05",  x"3e",  x"32", -- 1040
         x"32",  x"88",  x"00",  x"2b",  x"46",  x"2b",  x"4e",  x"30", -- 1048
         x"0d",  x"e1",  x"cd",  x"1a",  x"c9",  x"d5",  x"3e",  x"33", -- 1050
         x"32",  x"88",  x"00",  x"01",  x"00",  x"00",  x"21",  x"85", -- 1058
         x"00",  x"7e",  x"36",  x"00",  x"2a",  x"80",  x"00",  x"fe", -- 1060
         x"2d",  x"20",  x"04",  x"ed",  x"42",  x"18",  x"0a",  x"fe", -- 1068
         x"2b",  x"28",  x"05",  x"3e",  x"42",  x"32",  x"88",  x"00", -- 1070
         x"09",  x"22",  x"80",  x"00",  x"e1",  x"c3",  x"51",  x"cf", -- 1078
         x"d5",  x"c1",  x"18",  x"da",  x"f5",  x"23",  x"7e",  x"eb", -- 1080
         x"cd",  x"40",  x"c9",  x"30",  x"1b",  x"f1",  x"fe",  x"4d", -- 1088
         x"20",  x"08",  x"3e",  x"28",  x"32",  x"83",  x"00",  x"eb", -- 1090
         x"18",  x"5b",  x"21",  x"f9",  x"d0",  x"01",  x"09",  x"00", -- 1098
         x"ed",  x"b1",  x"20",  x"97",  x"cb",  x"21",  x"18",  x"20", -- 10A0
         x"13",  x"21",  x"08",  x"d1",  x"01",  x"0e",  x"00",  x"ed", -- 10A8
         x"b9",  x"20",  x"86",  x"d6",  x"19",  x"47",  x"cb",  x"41", -- 10B0
         x"ca",  x"39",  x"d0",  x"1a",  x"cd",  x"40",  x"c9",  x"d2", -- 10B8
         x"39",  x"d0",  x"f1",  x"be",  x"c2",  x"3a",  x"d0",  x"80", -- 10C0
         x"d6",  x"41",  x"06",  x"00",  x"eb",  x"32",  x"86",  x"00", -- 10C8
         x"fe",  x"3a",  x"20",  x"13",  x"3a",  x"83",  x"00",  x"b7", -- 10D0
         x"3e",  x"20",  x"28",  x"06",  x"af",  x"32",  x"83",  x"00", -- 10D8
         x"3e",  x"06",  x"32",  x"87",  x"00",  x"18",  x"96",  x"e5", -- 10E0
         x"21",  x"97",  x"d1",  x"09",  x"7e",  x"e1",  x"b7",  x"f2", -- 10E8
         x"e2",  x"d0",  x"32",  x"82",  x"00",  x"3e",  x"3a",  x"18", -- 10F0
         x"d4",  x"49",  x"52",  x"42",  x"43",  x"44",  x"45",  x"48", -- 10F8
         x"4c",  x"41",  x"46",  x"53",  x"50",  x"49",  x"58",  x"49", -- 1100
         x"59",  x"40",  x"b8",  x"40",  x"c2",  x"45",  x"38",  x"28", -- 1108
         x"18",  x"88",  x"80",  x"c4",  x"18",  x"05",  x"f4",  x"fc", -- 1110
         x"40",  x"00",  x"01",  x"70",  x"a0",  x"a9",  x"b9",  x"47", -- 1118
         x"aa",  x"98",  x"a1",  x"04",  x"ab",  x"a2",  x"00",  x"10", -- 1120
         x"30",  x"a3",  x"b0",  x"08",  x"68",  x"18",  x"20",  x"28", -- 1128
         x"08",  x"10",  x"77",  x"80",  x"c0",  x"c0",  x"01",  x"b2", -- 1130
         x"c1",  x"00",  x"38",  x"b3",  x"ba",  x"4e",  x"da",  x"10", -- 1138
         x"b1",  x"41",  x"46",  x"bb",  x"c8",  x"ac",  x"20",  x"b4", -- 1140
         x"bc",  x"c5",  x"a4",  x"a8",  x"00",  x"00",  x"02",  x"90", -- 1148
         x"43",  x"34",  x"76",  x"2a",  x"a3",  x"43",  x"33",  x"4c", -- 1150
         x"74",  x"04",  x"4a",  x"73",  x"54",  x"13",  x"33",  x"71", -- 1158
         x"42",  x"2d",  x"a3",  x"44",  x"c3",  x"e3",  x"f5",  x"83", -- 1160
         x"34",  x"93",  x"34",  x"c3",  x"d3",  x"29",  x"08",  x"03", -- 1168
         x"93",  x"04",  x"73",  x"83",  x"68",  x"53",  x"18",  x"78", -- 1170
         x"73",  x"03",  x"51",  x"6b",  x"21",  x"63",  x"c3",  x"63", -- 1178
         x"0f",  x"48",  x"c3",  x"93",  x"d3",  x"43",  x"6c",  x"b3", -- 1180
         x"27",  x"a3",  x"d3",  x"13",  x"83",  x"08",  x"c3",  x"93", -- 1188
         x"23",  x"d3",  x"14",  x"4e",  x"18",  x"6d",  x"24",  x"07", -- 1190
         x"00",  x"05",  x"10",  x"04",  x"20",  x"03",  x"30",  x"02", -- 1198
         x"30",  x"01",  x"dd",  x"00",  x"fd",  x"4f",  x"ff",  x"47", -- 11A0
         x"e2",  x"18",  x"16",  x"20",  x"8c",  x"7d",  x"58",  x"26", -- 11A8
         x"40",  x"4d",  x"61",  x"2e",  x"85",  x"63",  x"64",  x"8a", -- 11B0
         x"57",  x"98",  x"67",  x"72",  x"78",  x"94",  x"9a",  x"82", -- 11B8
         x"90",  x"24",  x"49",  x"65",  x"70",  x"3f",  x"00",  x"01", -- 11C0
         x"02",  x"03",  x"04",  x"05",  x"07",  x"0a",  x"43",  x"0b", -- 11C8
         x"0f",  x"3d",  x"44",  x"12",  x"15",  x"45",  x"23",  x"30", -- 11D0
         x"33",  x"46",  x"37",  x"3a",  x"3b",  x"42",  x"fe",  x"41", -- 11D8
         x"d8",  x"fe",  x"5b",  x"3f",  x"d0",  x"fe",  x"61",  x"d8", -- 11E0
         x"fe",  x"7b",  x"3f",  x"d8",  x"e6",  x"df",  x"c9",  x"06", -- 11E8
         x"01",  x"fe",  x"20",  x"30",  x"1c",  x"fe",  x"0d",  x"20", -- 11F0
         x"04",  x"16",  x"ff",  x"18",  x"14",  x"fe",  x"0a",  x"20", -- 11F8
         x"04",  x"15",  x"1c",  x"18",  x"0c",  x"fe",  x"09",  x"20", -- 1200
         x"06",  x"7a",  x"2f",  x"e6",  x"07",  x"3c",  x"47",  x"3e", -- 1208
         x"20",  x"c5",  x"d5",  x"e5",  x"cd",  x"03",  x"f0",  x"24", -- 1210
         x"e1",  x"d1",  x"c1",  x"14",  x"1d",  x"28",  x"02",  x"10", -- 1218
         x"f0",  x"cd",  x"03",  x"f0",  x"0c",  x"dd",  x"7e",  x"0d", -- 1220
         x"fe",  x"13",  x"c0",  x"c3",  x"63",  x"c7",  x"cd",  x"03", -- 1228
         x"f0",  x"20",  x"cd",  x"fe",  x"c5",  x"cd",  x"cb",  x"c5", -- 1230
         x"cd",  x"03",  x"f0",  x"23",  x"43",  x"4f",  x"4d",  x"00", -- 1238
         x"11",  x"00",  x"b7",  x"01",  x"0b",  x"00",  x"ed",  x"b0", -- 1240
         x"3e",  x"02",  x"32",  x"10",  x"b7",  x"2a",  x"7e",  x"00", -- 1248
         x"22",  x"13",  x"b7",  x"c9",  x"c5",  x"cb",  x"67",  x"28", -- 1250
         x"3f",  x"21",  x"00",  x"b7",  x"dd",  x"75",  x"05",  x"dd", -- 1258
         x"74",  x"06",  x"fd",  x"e5",  x"d1",  x"2a",  x"13",  x"b7", -- 1260
         x"19",  x"ed",  x"53",  x"11",  x"b7",  x"22",  x"13",  x"b7", -- 1268
         x"3e",  x"14",  x"32",  x"a0",  x"b7",  x"eb",  x"cd",  x"03", -- 1270
         x"f0",  x"1b",  x"cd",  x"03",  x"f0",  x"2c",  x"cd",  x"03", -- 1278
         x"f0",  x"08",  x"21",  x"6d",  x"00",  x"cb",  x"9e",  x"08", -- 1280
         x"af",  x"08",  x"dd",  x"7e",  x"02",  x"cd",  x"03",  x"f0", -- 1288
         x"1c",  x"cd",  x"03",  x"f0",  x"23",  x"20",  x"20",  x"00", -- 1290
         x"21",  x"00",  x"b7",  x"08",  x"fe",  x"80",  x"20",  x"09", -- 1298
         x"01",  x"a0",  x"00",  x"cd",  x"03",  x"f0",  x"01",  x"18", -- 12A0
         x"df",  x"6f",  x"3c",  x"08",  x"c1",  x"71",  x"c9",  x"fd", -- 12A8
         x"fd",  x"65",  x"01",  x"7d",  x"32",  x"f6",  x"b7",  x"c9", -- 12B0
         x"fd",  x"fd",  x"68",  x"01",  x"7d",  x"32",  x"f9",  x"b7", -- 12B8
         x"c9",  x"fd",  x"fd",  x"6c",  x"01",  x"7d",  x"32",  x"f8", -- 12C0
         x"b7",  x"c9",  x"fd",  x"fd",  x"62",  x"63",  x"01",  x"22", -- 12C8
         x"f4",  x"b7",  x"c9",  x"fd",  x"fd",  x"64",  x"65",  x"01", -- 12D0
         x"22",  x"f6",  x"b7",  x"c9",  x"fd",  x"fd",  x"68",  x"6c", -- 12D8
         x"01",  x"22",  x"f8",  x"b7",  x"c9",  x"fd",  x"fd",  x"69", -- 12E0
         x"79",  x"01",  x"e5",  x"fd",  x"e1",  x"c9",  x"fd",  x"fd", -- 12E8
         x"73",  x"70",  x"01",  x"22",  x"fc",  x"b7",  x"c9",  x"fd", -- 12F0
         x"fd",  x"70",  x"63",  x"01",  x"22",  x"fa",  x"b7",  x"c9", -- 12F8
         x"fd",  x"7e",  x"00",  x"fe",  x"dd",  x"20",  x"04",  x"1e", -- 1300
         x"80",  x"18",  x"06",  x"fe",  x"fd",  x"20",  x"0a",  x"1e", -- 1308
         x"c0",  x"fd",  x"7e",  x"02",  x"08",  x"fd",  x"23",  x"18", -- 1310
         x"e7",  x"21",  x"d2",  x"d3",  x"fe",  x"ed",  x"28",  x"13", -- 1318
         x"fe",  x"cb",  x"20",  x"18",  x"cb",  x"c3",  x"2e",  x"5a", -- 1320
         x"cb",  x"7b",  x"28",  x"0b",  x"fd",  x"23",  x"fd",  x"7e", -- 1328
         x"01",  x"18",  x"09",  x"2e",  x"7a",  x"1e",  x"20",  x"fd", -- 1330
         x"23",  x"fd",  x"7e",  x"00",  x"57",  x"cb",  x"7e",  x"23", -- 1338
         x"28",  x"fb",  x"7a",  x"ae",  x"23",  x"a6",  x"23",  x"20", -- 1340
         x"f4",  x"cd",  x"cf",  x"d4",  x"cd",  x"2a",  x"d5",  x"fd", -- 1348
         x"23",  x"d9",  x"c9",  x"4f",  x"d4",  x"7a",  x"0f",  x"0f", -- 1350
         x"0f",  x"a1",  x"c9",  x"00",  x"c0",  x"7b",  x"20",  x"f4", -- 1358
         x"40",  x"c0",  x"42",  x"49",  x"54",  x"20",  x"68",  x"2c", -- 1360
         x"f4",  x"80",  x"c0",  x"52",  x"45",  x"53",  x"20",  x"68", -- 1368
         x"2c",  x"f4",  x"c0",  x"c0",  x"53",  x"45",  x"54",  x"20", -- 1370
         x"68",  x"2c",  x"f4",  x"40",  x"c7",  x"1a",  x"66",  x"76", -- 1378
         x"0a",  x"43",  x"a9",  x"41",  x"c7",  x"1b",  x"66",  x"28", -- 1380
         x"43",  x"0b",  x"f6",  x"42",  x"cf",  x"1f",  x"66",  x"12", -- 1388
         x"2c",  x"eb",  x"4a",  x"cf",  x"1d",  x"66",  x"12",  x"2c", -- 1390
         x"eb",  x"4b",  x"cf",  x"01",  x"6b",  x"0a",  x"70",  x"a9", -- 1398
         x"43",  x"cf",  x"01",  x"28",  x"70",  x"0b",  x"eb",  x"44", -- 13A0
         x"c7",  x"4e",  x"45",  x"c7",  x"4d",  x"cf",  x"08",  x"49", -- 13A8
         x"a0",  x"45",  x"cf",  x"08",  x"4e",  x"a0",  x"46",  x"ff", -- 13B0
         x"0d",  x"b0",  x"56",  x"ff",  x"0d",  x"b1",  x"5e",  x"ff", -- 13B8
         x"0d",  x"b2",  x"47",  x"e7",  x"01",  x"f8",  x"67",  x"f7", -- 13C0
         x"77",  x"c4",  x"a0",  x"e4",  x"6a",  x"fa",  x"00",  x"00", -- 13C8
         x"3b",  x"66",  x"f2",  x"76",  x"ff",  x"48",  x"41",  x"4c", -- 13D0
         x"d4",  x"40",  x"c0",  x"01",  x"76",  x"2c",  x"f4",  x"06", -- 13D8
         x"c7",  x"01",  x"76",  x"2c",  x"ef",  x"02",  x"e7",  x"01", -- 13E0
         x"f9",  x"3a",  x"ff",  x"01",  x"41",  x"0a",  x"70",  x"a9", -- 13E8
         x"32",  x"ff",  x"01",  x"28",  x"70",  x"0b",  x"c1",  x"01", -- 13F0
         x"cf",  x"01",  x"6b",  x"2c",  x"f0",  x"2a",  x"ff",  x"01", -- 13F8
         x"75",  x"0a",  x"70",  x"a9",  x"22",  x"ff",  x"01",  x"28", -- 1400
         x"70",  x"0b",  x"f5",  x"f9",  x"ff",  x"01",  x"13",  x"2c", -- 1408
         x"f5",  x"f5",  x"ff",  x"05",  x"84",  x"c5",  x"cf",  x"05", -- 1410
         x"eb",  x"f1",  x"ff",  x"06",  x"84",  x"c1",  x"cf",  x"06", -- 1418
         x"eb",  x"20",  x"e7",  x"4a",  x"52",  x"66",  x"7e",  x"2c", -- 1420
         x"f1",  x"18",  x"ff",  x"4a",  x"52",  x"66",  x"71",  x"a0", -- 1428
         x"10",  x"ff",  x"44",  x"4a",  x"4e",  x"5a",  x"66",  x"f1", -- 1430
         x"cd",  x"ff",  x"07",  x"70",  x"a0",  x"c4",  x"c7",  x"07", -- 1438
         x"7d",  x"2c",  x"f0",  x"c9",  x"ff",  x"88",  x"c0",  x"c7", -- 1440
         x"08",  x"20",  x"7d",  x"e6",  x"e9",  x"ff",  x"0c",  x"6d", -- 1448
         x"a0",  x"04",  x"c6",  x"69",  x"f6",  x"09",  x"cf",  x"1c", -- 1450
         x"66",  x"75",  x"2c",  x"eb",  x"03",  x"cf",  x"16",  x"eb", -- 1458
         x"0b",  x"cf",  x"17",  x"eb",  x"80",  x"c0",  x"7f",  x"66", -- 1460
         x"f4",  x"c6",  x"c7",  x"7f",  x"66",  x"ef",  x"c3",  x"ff", -- 1468
         x"0c",  x"70",  x"a0",  x"c2",  x"c7",  x"0c",  x"7d",  x"2c", -- 1470
         x"f0",  x"eb",  x"ff",  x"09",  x"11",  x"2c",  x"92",  x"d9", -- 1478
         x"ff",  x"45",  x"58",  x"d8",  x"08",  x"ff",  x"09",  x"04", -- 1480
         x"2c",  x"04",  x"a7",  x"e3",  x"ff",  x"09",  x"28",  x"13", -- 1488
         x"0b",  x"f5",  x"07",  x"e7",  x"7c",  x"c1",  x"db",  x"ff", -- 1490
         x"1a",  x"66",  x"03",  x"ef",  x"d3",  x"ff",  x"1b",  x"66", -- 1498
         x"6f",  x"82",  x"27",  x"ff",  x"44",  x"41",  x"c1",  x"2f", -- 14A0
         x"ff",  x"19",  x"cc",  x"3f",  x"ff",  x"43",  x"43",  x"c6", -- 14A8
         x"f3",  x"ff",  x"44",  x"c9",  x"fb",  x"ff",  x"45",  x"c9", -- 14B0
         x"37",  x"ff",  x"53",  x"43",  x"c6",  x"c7",  x"c7",  x"52", -- 14B8
         x"53",  x"54",  x"66",  x"6c",  x"a0",  x"00",  x"ff",  x"4e", -- 14C0
         x"4f",  x"d0",  x"e1",  x"cb",  x"7e",  x"23",  x"c0",  x"7e", -- 14C8
         x"e5",  x"e6",  x"7f",  x"21",  x"ca",  x"d4",  x"e5",  x"fe", -- 14D0
         x"20",  x"38",  x"58",  x"fe",  x"60",  x"38",  x"52",  x"0e", -- 14D8
         x"07",  x"c6",  x"89",  x"38",  x"07",  x"21",  x"11",  x"d5", -- 14E0
         x"85",  x"6f",  x"6e",  x"e9",  x"21",  x"f4",  x"d6",  x"85", -- 14E8
         x"6f",  x"6e",  x"cd",  x"55",  x"d3",  x"3c",  x"cb",  x"7e", -- 14F0
         x"23",  x"28",  x"fb",  x"3d",  x"20",  x"f8",  x"18",  x"cf", -- 14F8
         x"25",  x"de",  x"11",  x"a4",  x"a9",  x"c2",  x"38",  x"4f", -- 1500
         x"51",  x"3d",  x"55",  x"6e",  x"16",  x"2a",  x"e0",  x"be", -- 1508
         x"db",  x"cd",  x"55",  x"d3",  x"18",  x"7c",  x"cb",  x"7b", -- 1510
         x"28",  x"06",  x"fd",  x"7e",  x"fe",  x"cd",  x"89",  x"d5", -- 1518
         x"6a",  x"26",  x"ed",  x"18",  x"5f",  x"3e",  x"20",  x"c3", -- 1520
         x"9a",  x"d5",  x"3e",  x"0d",  x"cd",  x"9a",  x"d5",  x"3e", -- 1528
         x"0a",  x"18",  x"67",  x"21",  x"50",  x"d6",  x"18",  x"bd", -- 1530
         x"7a",  x"e6",  x"38",  x"18",  x"0a",  x"fd",  x"23",  x"3e", -- 1538
         x"30",  x"cd",  x"9a",  x"d5",  x"fd",  x"7e",  x"00",  x"cd", -- 1540
         x"89",  x"d5",  x"3e",  x"48",  x"c3",  x"fe",  x"d6",  x"af", -- 1548
         x"08",  x"79",  x"c3",  x"e3",  x"d5",  x"fd",  x"23",  x"fd", -- 1550
         x"23",  x"fd",  x"66",  x"00",  x"fd",  x"6e",  x"ff",  x"3e", -- 1558
         x"30",  x"cd",  x"9a",  x"d5",  x"cd",  x"84",  x"d5",  x"18", -- 1560
         x"e1",  x"3e",  x"30",  x"cd",  x"9a",  x"d5",  x"fd",  x"23", -- 1568
         x"d9",  x"d5",  x"d9",  x"e1",  x"fd",  x"e5",  x"c1",  x"09", -- 1570
         x"23",  x"0a",  x"4f",  x"17",  x"06",  x"00",  x"30",  x"01", -- 1578
         x"05",  x"09",  x"18",  x"db",  x"7c",  x"cd",  x"89",  x"d5", -- 1580
         x"7d",  x"f5",  x"1f",  x"1f",  x"1f",  x"1f",  x"cd",  x"92", -- 1588
         x"d5",  x"f1",  x"e6",  x"0f",  x"c6",  x"90",  x"27",  x"ce", -- 1590
         x"40",  x"27",  x"e5",  x"d5",  x"c5",  x"cd",  x"fe",  x"d6", -- 1598
         x"c1",  x"d1",  x"e1",  x"c9",  x"21",  x"81",  x"d6",  x"18", -- 15A0
         x"0a",  x"21",  x"8f",  x"d6",  x"7a",  x"ee",  x"b3",  x"e6", -- 15A8
         x"f7",  x"28",  x"05",  x"7a",  x"a1",  x"c3",  x"36",  x"d5", -- 15B0
         x"21",  x"53",  x"d3",  x"c3",  x"cf",  x"d4",  x"3e",  x"02", -- 15B8
         x"18",  x"04",  x"cd",  x"55",  x"d3",  x"1f",  x"21",  x"7d", -- 15C0
         x"d6",  x"fe",  x"02",  x"20",  x"e8",  x"cb",  x"7b",  x"28", -- 15C8
         x"e4",  x"c6",  x"02",  x"cb",  x"73",  x"ca",  x"36",  x"d5", -- 15D0
         x"3c",  x"18",  x"da",  x"cd",  x"55",  x"d3",  x"18",  x"01", -- 15D8
         x"7a",  x"3c",  x"a1",  x"cb",  x"7b",  x"28",  x"27",  x"cb", -- 15E0
         x"43",  x"20",  x"50",  x"fe",  x"05",  x"38",  x"1f",  x"47", -- 15E8
         x"7a",  x"ee",  x"70",  x"e6",  x"78",  x"28",  x"3e",  x"7a", -- 15F0
         x"ee",  x"46",  x"e6",  x"c7",  x"28",  x"37",  x"78",  x"b9", -- 15F8
         x"20",  x"04",  x"cb",  x"cb",  x"fd",  x"23",  x"c6",  x"03", -- 1600
         x"cb",  x"73",  x"28",  x"02",  x"c6",  x"03",  x"21",  x"0b", -- 1608
         x"d7",  x"cd",  x"f5",  x"d4",  x"cb",  x"4b",  x"c8",  x"cb", -- 1610
         x"8b",  x"08",  x"b7",  x"28",  x"13",  x"47",  x"3e",  x"2b", -- 1618
         x"f2",  x"29",  x"d6",  x"78",  x"ed",  x"44",  x"47",  x"3e", -- 1620
         x"2d",  x"cd",  x"9a",  x"d5",  x"78",  x"cd",  x"47",  x"d5", -- 1628
         x"3e",  x"29",  x"c3",  x"9a",  x"d5",  x"78",  x"b9",  x"28", -- 1630
         x"c9",  x"18",  x"d3",  x"f5",  x"79",  x"cd",  x"02",  x"d6", -- 1638
         x"f1",  x"b9",  x"c8",  x"47",  x"7a",  x"ee",  x"40",  x"e6", -- 1640
         x"40",  x"c8",  x"af",  x"cd",  x"33",  x"d5",  x"78",  x"18", -- 1648
         x"bd",  x"26",  x"81",  x"18",  x"e6",  x"2c",  x"c1",  x"41", -- 1650
         x"ac",  x"41",  x"c6",  x"50",  x"55",  x"53",  x"48",  x"e6", -- 1658
         x"50",  x"4f",  x"50",  x"e6",  x"43",  x"41",  x"4c",  x"4c", -- 1660
         x"e6",  x"52",  x"45",  x"d4",  x"45",  x"58",  x"e6",  x"2c", -- 1668
         x"a8",  x"29",  x"ac",  x"4a",  x"50",  x"20",  x"e6",  x"49", -- 1670
         x"4d",  x"e6",  x"52",  x"d2",  x"52",  x"cc",  x"42",  x"c3", -- 1678
         x"44",  x"c5",  x"48",  x"cc",  x"53",  x"d0",  x"49",  x"d8", -- 1680
         x"49",  x"d9",  x"1a",  x"43",  x"e6",  x"11",  x"43",  x"e6", -- 1688
         x"4c",  x"c4",  x"43",  x"d0",  x"49",  x"ce",  x"4f",  x"55", -- 1690
         x"d4",  x"41",  x"44",  x"c4",  x"41",  x"44",  x"c3",  x"53", -- 1698
         x"55",  x"c2",  x"53",  x"90",  x"41",  x"4e",  x"c4",  x"58", -- 16A0
         x"4f",  x"d2",  x"4f",  x"d2",  x"43",  x"50",  x"a0",  x"fb", -- 16A8
         x"fb",  x"8f",  x"8e",  x"0f",  x"c3",  x"0e",  x"c3",  x"0f", -- 16B0
         x"a0",  x"0e",  x"a0",  x"53",  x"4c",  x"c1",  x"53",  x"52", -- 16B8
         x"c1",  x"53",  x"4c",  x"d3",  x"53",  x"8f",  x"c9",  x"c4", -- 16C0
         x"49",  x"d2",  x"44",  x"d2",  x"4e",  x"da",  x"da",  x"4e", -- 16C8
         x"c3",  x"c3",  x"50",  x"cf",  x"50",  x"c5",  x"d0",  x"cd", -- 16D0
         x"28",  x"10",  x"0b",  x"c1",  x"41",  x"0a",  x"10",  x"a9", -- 16D8
         x"28",  x"11",  x"0b",  x"c1",  x"41",  x"0a",  x"11",  x"a9", -- 16E0
         x"49",  x"2c",  x"c1",  x"52",  x"2c",  x"c1",  x"41",  x"2c", -- 16E8
         x"c9",  x"41",  x"2c",  x"d2",  x"6e",  x"e7",  x"d7",  x"ba", -- 16F0
         x"b2",  x"ae",  x"cb",  x"c5",  x"98",  x"00",  x"f5",  x"3a", -- 16F8
         x"fe",  x"b7",  x"a7",  x"c2",  x"21",  x"d8",  x"f1",  x"cd", -- 1700
         x"03",  x"f0",  x"24",  x"c9",  x"c1",  x"c2",  x"c3",  x"c4", -- 1708
         x"c5",  x"c8",  x"cc",  x"28",  x"12",  x"a9",  x"48",  x"d8", -- 1710
         x"4c",  x"d8",  x"28",  x"94",  x"48",  x"d9",  x"4c",  x"d9", -- 1718
         x"28",  x"95",  x"cd",  x"b6",  x"d7",  x"3e",  x"20",  x"cd", -- 1720
         x"9a",  x"d5",  x"3a",  x"ff",  x"b7",  x"a7",  x"20",  x"22", -- 1728
         x"fd",  x"e5",  x"e1",  x"06",  x"00",  x"7e",  x"fe",  x"cd", -- 1730
         x"20",  x"0e",  x"23",  x"7e",  x"fe",  x"03",  x"20",  x"08", -- 1738
         x"23",  x"7e",  x"fe",  x"f0",  x"20",  x"02",  x"06",  x"02", -- 1740
         x"78",  x"32",  x"ff",  x"b7",  x"d9",  x"1e",  x"00",  x"c3", -- 1748
         x"00",  x"d3",  x"3d",  x"28",  x"0e",  x"32",  x"ff",  x"b7", -- 1750
         x"cd",  x"9a",  x"d7",  x"fe",  x"23",  x"c8",  x"af",  x"32", -- 1758
         x"ff",  x"b7",  x"c9",  x"fd",  x"7e",  x"00",  x"fe",  x"20", -- 1760
         x"38",  x"29",  x"fe",  x"80",  x"30",  x"25",  x"21",  x"b1", -- 1768
         x"d7",  x"f5",  x"cd",  x"cf",  x"d4",  x"3e",  x"27",  x"cd", -- 1770
         x"fe",  x"d6",  x"f1",  x"cd",  x"fe",  x"d6",  x"fd",  x"23", -- 1778
         x"fd",  x"7e",  x"00",  x"fe",  x"20",  x"38",  x"04",  x"fe", -- 1780
         x"80",  x"38",  x"f0",  x"3e",  x"27",  x"cd",  x"fe",  x"d6", -- 1788
         x"c3",  x"2a",  x"d5",  x"cd",  x"9a",  x"d7",  x"a7",  x"c0", -- 1790
         x"18",  x"c4",  x"21",  x"ac",  x"d7",  x"cd",  x"cf",  x"d4", -- 1798
         x"cd",  x"3f",  x"d5",  x"cd",  x"2a",  x"d5",  x"fd",  x"7e", -- 17A0
         x"00",  x"fd",  x"23",  x"c9",  x"44",  x"45",  x"46",  x"42", -- 17A8
         x"a0",  x"44",  x"45",  x"46",  x"4d",  x"a0",  x"fd",  x"e5", -- 17B0
         x"e1",  x"19",  x"c3",  x"84",  x"d5",  x"7f",  x"7f",  x"44", -- 17B8
         x"49",  x"53",  x"41",  x"53",  x"53",  x"01",  x"af",  x"32", -- 17C0
         x"fe",  x"b7",  x"32",  x"ff",  x"b7",  x"e5",  x"fd",  x"e1", -- 17C8
         x"3a",  x"81",  x"b7",  x"fe",  x"03",  x"30",  x"07",  x"01", -- 17D0
         x"1c",  x"00",  x"ed",  x"43",  x"86",  x"b7",  x"fe",  x"04", -- 17D8
         x"11",  x"00",  x"00",  x"38",  x"04",  x"ed",  x"5b",  x"88", -- 17E0
         x"b7",  x"c5",  x"cd",  x"22",  x"d7",  x"fd",  x"e5",  x"e1", -- 17E8
         x"ed",  x"5b",  x"84",  x"b7",  x"c1",  x"a7",  x"ed",  x"52", -- 17F0
         x"d0",  x"cd",  x"03",  x"f0",  x"2a",  x"d8",  x"0d",  x"3a", -- 17F8
         x"81",  x"b7",  x"c2",  x"de",  x"d7",  x"cd",  x"03",  x"f0", -- 1800
         x"04",  x"fe",  x"03",  x"c8",  x"fe",  x"0c",  x"20",  x"06", -- 1808
         x"cd",  x"03",  x"f0",  x"24",  x"18",  x"04",  x"fe",  x"0d", -- 1810
         x"20",  x"eb",  x"ed",  x"4b",  x"86",  x"b7",  x"c3",  x"d0", -- 1818
         x"d7",  x"f1",  x"2a",  x"97",  x"b7",  x"77",  x"3a",  x"96", -- 1820
         x"b7",  x"3d",  x"23",  x"20",  x"0c",  x"01",  x"e8",  x"03", -- 1828
         x"cd",  x"03",  x"f0",  x"01",  x"21",  x"00",  x"b7",  x"3e", -- 1830
         x"80",  x"22",  x"97",  x"b7",  x"32",  x"96",  x"b7",  x"c9", -- 1838
         x"7f",  x"7f",  x"43",  x"44",  x"49",  x"53",  x"41",  x"53", -- 1840
         x"53",  x"01",  x"e5",  x"fd",  x"e1",  x"cd",  x"03",  x"f0", -- 1848
         x"23",  x"4e",  x"41",  x"4d",  x"45",  x"20",  x"3a",  x"20", -- 1850
         x"00",  x"cd",  x"03",  x"f0",  x"17",  x"21",  x"07",  x"00", -- 1858
         x"19",  x"11",  x"00",  x"b7",  x"01",  x"08",  x"00",  x"ed", -- 1860
         x"b0",  x"eb",  x"36",  x"41",  x"23",  x"36",  x"53",  x"23", -- 1868
         x"36",  x"4d",  x"23",  x"af",  x"77",  x"32",  x"10",  x"b7", -- 1870
         x"32",  x"ff",  x"b7",  x"3c",  x"32",  x"fe",  x"b7",  x"cd", -- 1878
         x"03",  x"f0",  x"08",  x"cd",  x"34",  x"d8",  x"cd",  x"2a", -- 1880
         x"d5",  x"ed",  x"5b",  x"86",  x"b7",  x"3e",  x"09",  x"cd", -- 1888
         x"27",  x"d7",  x"fd",  x"e5",  x"e1",  x"ed",  x"4b",  x"84", -- 1890
         x"b7",  x"ed",  x"42",  x"38",  x"ec",  x"3e",  x"20",  x"cd", -- 1898
         x"9a",  x"d5",  x"3e",  x"03",  x"cd",  x"9a",  x"d5",  x"01", -- 18A0
         x"e8",  x"03",  x"cd",  x"03",  x"f0",  x"09",  x"c9",  x"06", -- 18A8
         x"04",  x"7e",  x"fe",  x"ed",  x"28",  x"2e",  x"cb",  x"af", -- 18B0
         x"fe",  x"dd",  x"28",  x"09",  x"7e",  x"fe",  x"cb",  x"20", -- 18B8
         x"2f",  x"06",  x"02",  x"18",  x"53",  x"23",  x"7e",  x"fe", -- 18C0
         x"cb",  x"28",  x"4d",  x"04",  x"e6",  x"f8",  x"fe",  x"30", -- 18C8
         x"28",  x"20",  x"fe",  x"70",  x"28",  x"1c",  x"7e",  x"e6", -- 18D0
         x"c7",  x"fe",  x"46",  x"28",  x"15",  x"fe",  x"86",  x"28", -- 18D8
         x"11",  x"05",  x"18",  x"0e",  x"23",  x"7e",  x"e6",  x"c7", -- 18E0
         x"fe",  x"43",  x"28",  x"2c",  x"06",  x"02",  x"18",  x"28", -- 18E8
         x"06",  x"03",  x"7e",  x"fe",  x"cd",  x"28",  x"1f",  x"fe", -- 18F0
         x"c3",  x"28",  x"1b",  x"e6",  x"e7",  x"fe",  x"22",  x"28", -- 18F8
         x"17",  x"7e",  x"e6",  x"cf",  x"fe",  x"01",  x"28",  x"10", -- 1900
         x"05",  x"e6",  x"c7",  x"28",  x"20",  x"fe",  x"c2",  x"28", -- 1908
         x"04",  x"fe",  x"c4",  x"20",  x"05",  x"04",  x"af",  x"c9", -- 1910
         x"a7",  x"c9",  x"fe",  x"06",  x"28",  x"fa",  x"fe",  x"c6", -- 1918
         x"28",  x"f6",  x"7e",  x"e6",  x"f7",  x"fe",  x"d3",  x"28", -- 1920
         x"ef",  x"05",  x"78",  x"18",  x"eb",  x"7e",  x"fe",  x"09", -- 1928
         x"38",  x"f7",  x"37",  x"c9",  x"fd",  x"fd",  x"4d",  x"45", -- 1930
         x"4e",  x"55",  x"01",  x"e1",  x"18",  x"38",  x"7f",  x"7f", -- 1938
         x"54",  x"45",  x"4d",  x"4f",  x"01",  x"3a",  x"81",  x"b7", -- 1940
         x"a7",  x"3e",  x"ff",  x"20",  x"01",  x"af",  x"32",  x"ed", -- 1948
         x"b7",  x"21",  x"ee",  x"b7",  x"06",  x"10",  x"36",  x"00", -- 1950
         x"23",  x"10",  x"fb",  x"2e",  x"60",  x"3a",  x"d7",  x"b7", -- 1958
         x"67",  x"22",  x"fc",  x"b7",  x"18",  x"09",  x"7f",  x"7f", -- 1960
         x"52",  x"45",  x"54",  x"45",  x"4d",  x"4f",  x"01",  x"2e", -- 1968
         x"e8",  x"36",  x"16",  x"23",  x"36",  x"da",  x"cd",  x"03", -- 1970
         x"f0",  x"23",  x"0c",  x"20",  x"3e",  x"3e",  x"3e",  x"20", -- 1978
         x"54",  x"45",  x"4d",  x"4f",  x"20",  x"3c",  x"3c",  x"3c", -- 1980
         x"00",  x"3a",  x"ed",  x"b7",  x"a7",  x"20",  x"0f",  x"cd", -- 1988
         x"03",  x"f0",  x"23",  x"20",  x"20",  x"28",  x"44",  x"49", -- 1990
         x"53",  x"41",  x"53",  x"53",  x"29",  x"00",  x"cd",  x"03", -- 1998
         x"f0",  x"2c",  x"21",  x"00",  x"ba",  x"01",  x"00",  x"26", -- 19A0
         x"cd",  x"03",  x"f0",  x"23",  x"0d",  x"02",  x"2b",  x"00", -- 19A8
         x"cd",  x"03",  x"f0",  x"2a",  x"38",  x"2c",  x"3e",  x"fd", -- 19B0
         x"ed",  x"b1",  x"e2",  x"e2",  x"d9",  x"ed",  x"a1",  x"20", -- 19B8
         x"f7",  x"7e",  x"fe",  x"02",  x"38",  x"10",  x"fe",  x"30", -- 19C0
         x"38",  x"de",  x"fe",  x"5f",  x"30",  x"da",  x"cd",  x"03", -- 19C8
         x"f0",  x"24",  x"23",  x"0b",  x"18",  x"eb",  x"cd",  x"03", -- 19D0
         x"f0",  x"2c",  x"18",  x"cc",  x"cd",  x"03",  x"f0",  x"23", -- 19D8
         x"2b",  x"00",  x"cd",  x"03",  x"f0",  x"17",  x"13",  x"1a", -- 19E0
         x"fe",  x"20",  x"28",  x"f0",  x"a7",  x"28",  x"ed",  x"3e", -- 19E8
         x"fd",  x"21",  x"00",  x"ba",  x"01",  x"00",  x"26",  x"cd", -- 19F0
         x"03",  x"f0",  x"1d",  x"30",  x"08",  x"e5",  x"cd",  x"03", -- 19F8
         x"f0",  x"22",  x"30",  x"07",  x"e1",  x"cd",  x"03",  x"f0", -- 1A00
         x"19",  x"18",  x"d1",  x"21",  x"dc",  x"d9",  x"e3",  x"23", -- 1A08
         x"e5",  x"cd",  x"03",  x"f0",  x"15",  x"c9",  x"e5",  x"21", -- 1A10
         x"27",  x"da",  x"e3",  x"f5",  x"3e",  x"03",  x"d3",  x"8c", -- 1A18
         x"f1",  x"fb",  x"ed",  x"4d",  x"e3",  x"2b",  x"e3",  x"22", -- 1A20
         x"f8",  x"b7",  x"f5",  x"e1",  x"22",  x"f2",  x"b7",  x"ed", -- 1A28
         x"53",  x"f6",  x"b7",  x"ed",  x"43",  x"f4",  x"b7",  x"e1", -- 1A30
         x"22",  x"fa",  x"b7",  x"21",  x"00",  x"00",  x"39",  x"22", -- 1A38
         x"fc",  x"b7",  x"ed",  x"7b",  x"ae",  x"b7",  x"3a",  x"ea", -- 1A40
         x"b7",  x"a7",  x"28",  x"16",  x"cd",  x"03",  x"f0",  x"2a", -- 1A48
         x"38",  x"0c",  x"2a",  x"fa",  x"b7",  x"ed",  x"5b",  x"eb", -- 1A50
         x"b7",  x"ed",  x"52",  x"c2",  x"0a",  x"dc",  x"af",  x"32", -- 1A58
         x"ea",  x"b7",  x"06",  x"06",  x"21",  x"f2",  x"b7",  x"cd", -- 1A60
         x"03",  x"f0",  x"23",  x"20",  x"41",  x"46",  x"20",  x"20", -- 1A68
         x"20",  x"42",  x"43",  x"20",  x"20",  x"20",  x"44",  x"45", -- 1A70
         x"20",  x"20",  x"20",  x"48",  x"4c",  x"20",  x"20",  x"20", -- 1A78
         x"50",  x"43",  x"20",  x"20",  x"20",  x"53",  x"50",  x"20", -- 1A80
         x"20",  x"20",  x"49",  x"0d",  x"0a",  x"00",  x"5e",  x"23", -- 1A88
         x"56",  x"23",  x"eb",  x"cd",  x"03",  x"f0",  x"1a",  x"eb", -- 1A90
         x"10",  x"f4",  x"ed",  x"57",  x"cd",  x"03",  x"f0",  x"1c", -- 1A98
         x"cd",  x"03",  x"f0",  x"2c",  x"cd",  x"03",  x"f0",  x"23", -- 1AA0
         x"20",  x"49",  x"58",  x"20",  x"20",  x"20",  x"49",  x"59", -- 1AA8
         x"20",  x"46",  x"4c",  x"41",  x"47",  x"53",  x"20",  x"4f", -- 1AB0
         x"50",  x"2e",  x"43",  x"4f",  x"44",  x"45",  x"0d",  x"0a", -- 1AB8
         x"00",  x"dd",  x"e5",  x"e1",  x"cd",  x"03",  x"f0",  x"1a", -- 1AC0
         x"fd",  x"e5",  x"e1",  x"cd",  x"03",  x"f0",  x"1a",  x"3a", -- 1AC8
         x"f2",  x"b7",  x"11",  x"76",  x"db",  x"06",  x"08",  x"13", -- 1AD0
         x"17",  x"f5",  x"1a",  x"30",  x"04",  x"cd",  x"03",  x"f0", -- 1AD8
         x"24",  x"f1",  x"10",  x"f3",  x"cd",  x"03",  x"f0",  x"23", -- 1AE0
         x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"00",  x"3a", -- 1AE8
         x"f1",  x"b7",  x"a7",  x"c4",  x"dd",  x"db",  x"af",  x"32", -- 1AF0
         x"f1",  x"b7",  x"2a",  x"fa",  x"b7",  x"e5",  x"cd",  x"af", -- 1AF8
         x"d8",  x"e1",  x"7e",  x"cd",  x"03",  x"f0",  x"1c",  x"23", -- 1B00
         x"10",  x"f8",  x"cd",  x"03",  x"f0",  x"2c",  x"3a",  x"ed", -- 1B08
         x"b7",  x"a7",  x"20",  x"12",  x"fd",  x"e5",  x"fd",  x"2a", -- 1B10
         x"fa",  x"b7",  x"11",  x"00",  x"00",  x"af",  x"32",  x"ff", -- 1B18
         x"b7",  x"cd",  x"22",  x"d7",  x"fd",  x"e1",  x"cd",  x"03", -- 1B20
         x"f0",  x"04",  x"fe",  x"0d",  x"ca",  x"74",  x"db",  x"fe", -- 1B28
         x"0a",  x"28",  x"07",  x"fe",  x"03",  x"20",  x"ef",  x"c3", -- 1B30
         x"dc",  x"d9",  x"3e",  x"01",  x"32",  x"ea",  x"b7",  x"2a", -- 1B38
         x"fa",  x"b7",  x"e5",  x"7e",  x"fe",  x"cd",  x"20",  x"1c", -- 1B40
         x"23",  x"7e",  x"fe",  x"03",  x"20",  x"16",  x"23",  x"7e", -- 1B48
         x"fe",  x"f0",  x"20",  x"10",  x"06",  x"04",  x"23",  x"7e", -- 1B50
         x"fe",  x"23",  x"20",  x"0d",  x"04",  x"23",  x"7e",  x"a7", -- 1B58
         x"20",  x"fa",  x"18",  x"05",  x"e1",  x"e5",  x"cd",  x"af", -- 1B60
         x"d8",  x"e1",  x"7d",  x"80",  x"6f",  x"3e",  x"00",  x"8c", -- 1B68
         x"67",  x"22",  x"eb",  x"b7",  x"c3",  x"0a",  x"dc",  x"53", -- 1B70
         x"5a",  x"00",  x"48",  x"00",  x"50",  x"4e",  x"43",  x"fd", -- 1B78
         x"fd",  x"41",  x"52",  x"49",  x"54",  x"48",  x"01",  x"eb", -- 1B80
         x"e5",  x"19",  x"cd",  x"03",  x"f0",  x"1a",  x"e1",  x"b7", -- 1B88
         x"ed",  x"52",  x"cd",  x"03",  x"f0",  x"1a",  x"2b",  x"2b", -- 1B90
         x"7c",  x"fe",  x"ff",  x"20",  x"0e",  x"cb",  x"7d",  x"20", -- 1B98
         x"11",  x"cd",  x"03",  x"f0",  x"23",  x"3f",  x"3f",  x"0d", -- 1BA0
         x"0a",  x"00",  x"c9",  x"b7",  x"20",  x"f3",  x"cb",  x"7d", -- 1BA8
         x"20",  x"ef",  x"7d",  x"cd",  x"03",  x"f0",  x"1c",  x"cd", -- 1BB0
         x"03",  x"f0",  x"2c",  x"c9",  x"fd",  x"fd",  x"42",  x"52", -- 1BB8
         x"45",  x"41",  x"4b",  x"01",  x"22",  x"ee",  x"b7",  x"3e", -- 1BC0
         x"c3",  x"21",  x"24",  x"da",  x"32",  x"38",  x"00",  x"22", -- 1BC8
         x"39",  x"00",  x"c9",  x"2a",  x"ee",  x"b7",  x"7e",  x"32", -- 1BD0
         x"f0",  x"b7",  x"36",  x"ff",  x"c9",  x"2a",  x"ee",  x"b7", -- 1BD8
         x"3a",  x"f0",  x"b7",  x"77",  x"c9",  x"fd",  x"fd",  x"47", -- 1BE0
         x"4f",  x"01",  x"3e",  x"ff",  x"32",  x"f1",  x"b7",  x"e5", -- 1BE8
         x"cd",  x"d3",  x"db",  x"e1",  x"18",  x"0b",  x"fd",  x"fd", -- 1BF0
         x"53",  x"54",  x"45",  x"50",  x"01",  x"af",  x"32",  x"f1", -- 1BF8
         x"b7",  x"3a",  x"81",  x"b7",  x"b7",  x"28",  x"03",  x"22", -- 1C00
         x"fa",  x"b7",  x"ed",  x"4b",  x"f4",  x"b7",  x"ed",  x"5b", -- 1C08
         x"f6",  x"b7",  x"2a",  x"f2",  x"b7",  x"e5",  x"f1",  x"2a", -- 1C10
         x"fc",  x"b7",  x"f9",  x"2a",  x"fa",  x"b7",  x"e5",  x"2a", -- 1C18
         x"f8",  x"b7",  x"f5",  x"3a",  x"f1",  x"b7",  x"a7",  x"20", -- 1C20
         x"09",  x"3e",  x"87",  x"d3",  x"8c",  x"3e",  x"02",  x"d3", -- 1C28
         x"8c",  x"00",  x"f1",  x"00",  x"00",  x"c9",  x"fd",  x"fd", -- 1C30
         x"43",  x"4f",  x"50",  x"59",  x"01",  x"ed",  x"b0",  x"c9", -- 1C38
         x"fd",  x"fd",  x"4d",  x"4f",  x"56",  x"45",  x"01",  x"a7", -- 1C40
         x"ed",  x"52",  x"19",  x"30",  x"f0",  x"0b",  x"eb",  x"09", -- 1C48
         x"eb",  x"09",  x"03",  x"ed",  x"b8",  x"c9",  x"fd",  x"fd", -- 1C50
         x"52",  x"45",  x"47",  x"01",  x"7d",  x"fe",  x"06",  x"28", -- 1C58
         x"07",  x"38",  x"09",  x"cd",  x"03",  x"f0",  x"19",  x"c9", -- 1C60
         x"d5",  x"fd",  x"e1",  x"c9",  x"a7",  x"17",  x"21",  x"f2", -- 1C68
         x"b7",  x"85",  x"6f",  x"73",  x"23",  x"72",  x"c9",  x"fd", -- 1C70
         x"fd",  x"53",  x"42",  x"52",  x"4b",  x"01",  x"3e",  x"01", -- 1C78
         x"32",  x"ea",  x"b7",  x"22",  x"eb",  x"b7",  x"c9",  x"fd", -- 1C80
         x"fd",  x"49",  x"4e",  x"01",  x"e5",  x"c1",  x"ed",  x"78", -- 1C88
         x"cd",  x"03",  x"f0",  x"1c",  x"cd",  x"03",  x"f0",  x"2c", -- 1C90
         x"c9",  x"fd",  x"fd",  x"4f",  x"55",  x"54",  x"01",  x"e5", -- 1C98
         x"c1",  x"ed",  x"59",  x"c9",  x"fd",  x"fd",  x"44",  x"49", -- 1CA0
         x"53",  x"50",  x"4c",  x"41",  x"59",  x"01",  x"3a",  x"81", -- 1CA8
         x"b7",  x"fe",  x"03",  x"30",  x"02",  x"0e",  x"08",  x"c5", -- 1CB0
         x"cd",  x"03",  x"f0",  x"1a",  x"3e",  x"bf",  x"bc",  x"38", -- 1CB8
         x"4f",  x"e5",  x"06",  x"08",  x"7e",  x"cd",  x"03",  x"f0", -- 1CC0
         x"1c",  x"05",  x"28",  x"07",  x"cd",  x"03",  x"f0",  x"2b", -- 1CC8
         x"23",  x"18",  x"f1",  x"3e",  x"09",  x"cd",  x"03",  x"f0", -- 1CD0
         x"24",  x"cd",  x"f3",  x"dd",  x"e1",  x"06",  x"08",  x"7e", -- 1CD8
         x"cd",  x"03",  x"f0",  x"24",  x"23",  x"10",  x"f8",  x"cd", -- 1CE0
         x"f3",  x"dd",  x"cd",  x"03",  x"f0",  x"2c",  x"cd",  x"03", -- 1CE8
         x"f0",  x"2a",  x"38",  x"1c",  x"d5",  x"eb",  x"ed",  x"52", -- 1CF0
         x"eb",  x"d1",  x"38",  x"14",  x"0d",  x"20",  x"b9",  x"cd", -- 1CF8
         x"03",  x"f0",  x"04",  x"fe",  x"03",  x"c1",  x"c8",  x"fe", -- 1D00
         x"13",  x"20",  x"ac",  x"cd",  x"03",  x"f0",  x"2e",  x"c9", -- 1D08
         x"c1",  x"c9",  x"fd",  x"fd",  x"45",  x"58",  x"49",  x"54", -- 1D10
         x"01",  x"f1",  x"cd",  x"03",  x"f0",  x"12",  x"fd",  x"fd", -- 1D18
         x"4d",  x"4f",  x"44",  x"49",  x"46",  x"59",  x"01",  x"cd", -- 1D20
         x"03",  x"f0",  x"2e",  x"c9",  x"dd",  x"dd",  x"56",  x"45", -- 1D28
         x"52",  x"49",  x"46",  x"59",  x"01",  x"cd",  x"03",  x"f0", -- 1D30
         x"11",  x"c9",  x"fd",  x"fd",  x"46",  x"49",  x"4c",  x"4c", -- 1D38
         x"01",  x"eb",  x"a7",  x"ed",  x"52",  x"d8",  x"eb",  x"7b", -- 1D40
         x"b2",  x"c8",  x"71",  x"23",  x"1b",  x"18",  x"f8",  x"fd", -- 1D48
         x"fd",  x"43",  x"48",  x"53",  x"55",  x"4d",  x"01",  x"d5", -- 1D50
         x"c1",  x"cd",  x"83",  x"dd",  x"eb",  x"cd",  x"03",  x"f0", -- 1D58
         x"1a",  x"c3",  x"94",  x"dc",  x"fd",  x"fd",  x"57",  x"4f", -- 1D60
         x"52",  x"4b",  x"52",  x"41",  x"4d",  x"01",  x"f3",  x"65", -- 1D68
         x"7d",  x"32",  x"d7",  x"b7",  x"2e",  x"d4",  x"f9",  x"22", -- 1D70
         x"ae",  x"b7",  x"7c",  x"cd",  x"03",  x"f0",  x"31",  x"fb", -- 1D78
         x"c3",  x"5b",  x"d9",  x"11",  x"ff",  x"ff",  x"7e",  x"aa", -- 1D80
         x"57",  x"0f",  x"0f",  x"0f",  x"0f",  x"e6",  x"0f",  x"aa", -- 1D88
         x"57",  x"0f",  x"0f",  x"0f",  x"f5",  x"e6",  x"1f",  x"ab", -- 1D90
         x"5f",  x"f1",  x"f5",  x"0f",  x"e6",  x"f0",  x"ab",  x"5f", -- 1D98
         x"f1",  x"e6",  x"e0",  x"aa",  x"53",  x"5f",  x"23",  x"0b", -- 1DA0
         x"78",  x"b1",  x"20",  x"da",  x"c9",  x"fd",  x"fd",  x"63", -- 1DA8
         x"79",  x"01",  x"3a",  x"f2",  x"b7",  x"cb",  x"87",  x"06", -- 1DB0
         x"01",  x"cb",  x"45",  x"28",  x"01",  x"b0",  x"32",  x"f2", -- 1DB8
         x"b7",  x"c9",  x"fd",  x"fd",  x"7a",  x"01",  x"3a",  x"f2", -- 1DC0
         x"b7",  x"cb",  x"b7",  x"06",  x"40",  x"18",  x"ea",  x"fd", -- 1DC8
         x"fd",  x"61",  x"01",  x"7d",  x"32",  x"f3",  x"b7",  x"c9", -- 1DD0
         x"fd",  x"fd",  x"62",  x"01",  x"7d",  x"32",  x"f5",  x"b7", -- 1DD8
         x"c9",  x"fd",  x"fd",  x"63",  x"01",  x"7d",  x"32",  x"f4", -- 1DE0
         x"b7",  x"c9",  x"fd",  x"fd",  x"64",  x"01",  x"7d",  x"32", -- 1DE8
         x"f7",  x"b7",  x"c9",  x"f5",  x"3a",  x"a2",  x"b7",  x"ee", -- 1DF0
         x"08",  x"32",  x"a2",  x"b7",  x"f1",  x"c9",  x"ff",  x"ff", -- 1DF8
         x"07",  x"59",  x"04",  x"04",  x"03",  x"20",  x"05",  x"6a", -- 1E00
         x"1b",  x"5b",  x"31",  x"34",  x"34",  x"7d",  x"1b",  x"5b", -- 1E08
         x"31",  x"33",  x"32",  x"7a",  x"1b",  x"5b",  x"31",  x"32", -- 1E10
         x"60",  x"47",  x"5b",  x"04",  x"04",  x"03",  x"20",  x"05", -- 1E18
         x"6a",  x"7f",  x"7f",  x"56",  x"32",  x"34",  x"4b",  x"36", -- 1E20
         x"33",  x"31",  x"31",  x"01",  x"06",  x"11",  x"c5",  x"21", -- 1E28
         x"08",  x"de",  x"e5",  x"21",  x"00",  x"de",  x"e5",  x"18", -- 1E30
         x"16",  x"7f",  x"7f",  x"56",  x"32",  x"34",  x"4b",  x"36", -- 1E38
         x"33",  x"31",  x"33",  x"01",  x"06",  x"05",  x"c5",  x"21", -- 1E40
         x"13",  x"df",  x"e5",  x"21",  x"19",  x"de",  x"e5",  x"01", -- 1E48
         x"80",  x"08",  x"ed",  x"78",  x"fe",  x"ee",  x"28",  x"12", -- 1E50
         x"fe",  x"ff",  x"20",  x"08",  x"cd",  x"03",  x"f0",  x"19", -- 1E58
         x"e1",  x"e1",  x"e1",  x"c9",  x"3e",  x"04",  x"80",  x"47", -- 1E60
         x"18",  x"e8",  x"68",  x"3e",  x"02",  x"16",  x"01",  x"5a", -- 1E68
         x"cd",  x"03",  x"f0",  x"26",  x"cd",  x"95",  x"de",  x"21", -- 1E70
         x"a3",  x"de",  x"22",  x"99",  x"b7",  x"0e",  x"0c",  x"06", -- 1E78
         x"02",  x"e1",  x"f3",  x"ed",  x"b3",  x"01",  x"0a",  x"06", -- 1E80
         x"ed",  x"b3",  x"fb",  x"e1",  x"c1",  x"7e",  x"23",  x"cd", -- 1E88
         x"f7",  x"de",  x"10",  x"f9",  x"c9",  x"21",  x"c2",  x"de", -- 1E90
         x"11",  x"c4",  x"de",  x"22",  x"b9",  x"b7",  x"ed",  x"53", -- 1E98
         x"be",  x"b7",  x"c9",  x"e5",  x"d5",  x"2a",  x"b9",  x"b7", -- 1EA0
         x"6e",  x"2c",  x"2d",  x"20",  x"0c",  x"11",  x"be",  x"de", -- 1EA8
         x"21",  x"6c",  x"de",  x"cd",  x"9b",  x"de",  x"d1",  x"e1", -- 1EB0
         x"c9",  x"cd",  x"95",  x"de",  x"18",  x"f8",  x"f5",  x"cd", -- 1EB8
         x"03",  x"f0",  x"00",  x"f1",  x"f5",  x"3a",  x"a2",  x"b7", -- 1EC0
         x"cb",  x"5f",  x"28",  x"11",  x"f1",  x"f5",  x"fe",  x"7e", -- 1EC8
         x"30",  x"04",  x"fe",  x"20",  x"30",  x"22",  x"3e",  x"5f", -- 1ED0
         x"cd",  x"f7",  x"de",  x"f1",  x"c9",  x"f1",  x"fe",  x"0d", -- 1ED8
         x"20",  x"0f",  x"f5",  x"cd",  x"f7",  x"de",  x"3e",  x"20", -- 1EE0
         x"06",  x"0a",  x"cd",  x"f7",  x"de",  x"10",  x"fb",  x"18", -- 1EE8
         x"e7",  x"fe",  x"09",  x"20",  x"02",  x"3e",  x"20",  x"f5", -- 1EF0
         x"c5",  x"0e",  x"0a",  x"ed",  x"78",  x"cb",  x"57",  x"20", -- 1EF8
         x"09",  x"3e",  x"01",  x"cd",  x"03",  x"f0",  x"14",  x"c1", -- 1F00
         x"18",  x"ee",  x"c1",  x"f1",  x"c5",  x"0e",  x"08",  x"ed", -- 1F08
         x"79",  x"c1",  x"c9",  x"0d",  x"09",  x"1b",  x"4a",  x"18", -- 1F10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FF0
         x"d7",  x"61",  x"1c",  x"46",  x"39",  x"3d",  x"86",  x"07"  -- 1FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
