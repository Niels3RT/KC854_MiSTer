library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity caos47_e is
    generic(
        ADDR_WIDTH   : integer := 13
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end caos47_e;

architecture rtl of caos47_e is
    type rom8192x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom8192x8 := (
         x"c3",  x"66",  x"f1",  x"c3",  x"b6",  x"e5",  x"c3",  x"d3", -- 0000
         x"e5",  x"c3",  x"ba",  x"eb",  x"cf",  x"fc",  x"c3",  x"8a", -- 0008
         x"f8",  x"7f",  x"7f",  x"42",  x"41",  x"53",  x"49",  x"43", -- 0010
         x"11",  x"cd",  x"2f",  x"e0",  x"c3",  x"0d",  x"c0",  x"7f", -- 0018
         x"7f",  x"52",  x"45",  x"42",  x"41",  x"53",  x"49",  x"43", -- 0020
         x"11",  x"cd",  x"2f",  x"e0",  x"c3",  x"8c",  x"c0",  x"16", -- 0028
         x"00",  x"2e",  x"05",  x"cd",  x"02",  x"f1",  x"16",  x"c1", -- 0030
         x"cd",  x"00",  x"f1",  x"c3",  x"3f",  x"f0",  x"ed",  x"5b", -- 0038
         x"a0",  x"b7",  x"2a",  x"9c",  x"b7",  x"19",  x"cb",  x"24", -- 0040
         x"cb",  x"24",  x"cb",  x"24",  x"f5",  x"7d",  x"6c",  x"fe", -- 0048
         x"28",  x"30",  x"06",  x"f6",  x"80",  x"67",  x"f1",  x"a7", -- 0050
         x"c9",  x"f1",  x"37",  x"c9",  x"3a",  x"9e",  x"b7",  x"3d", -- 0058
         x"93",  x"d8",  x"3a",  x"9f",  x"b7",  x"3d",  x"92",  x"c9", -- 0060
         x"f5",  x"cd",  x"5c",  x"e0",  x"38",  x"eb",  x"3a",  x"9c", -- 0068
         x"b7",  x"83",  x"d5",  x"5f",  x"3a",  x"9d",  x"b7",  x"82", -- 0070
         x"87",  x"87",  x"87",  x"6f",  x"26",  x"00",  x"54",  x"29", -- 0078
         x"29",  x"19",  x"5f",  x"3a",  x"cc",  x"b7",  x"57",  x"19", -- 0080
         x"d1",  x"f1",  x"a7",  x"c9",  x"e5",  x"d5",  x"c5",  x"f5", -- 0088
         x"cd",  x"78",  x"e1",  x"ed",  x"53",  x"a0",  x"b7",  x"f1", -- 0090
         x"c1",  x"d1",  x"e1",  x"c9",  x"e5",  x"d5",  x"c5",  x"f5", -- 0098
         x"4f",  x"2a",  x"9c",  x"b7",  x"19",  x"eb",  x"7b",  x"fe", -- 00A0
         x"28",  x"30",  x"ec",  x"21",  x"a2",  x"b7",  x"cb",  x"6e", -- 00A8
         x"20",  x"63",  x"79",  x"21",  x"a6",  x"b7",  x"87",  x"30", -- 00B0
         x"02",  x"2e",  x"aa",  x"d6",  x"40",  x"f2",  x"c4",  x"e0", -- 00B8
         x"2c",  x"2c",  x"ee",  x"c0",  x"4e",  x"2c",  x"46",  x"87", -- 00C0
         x"6f",  x"26",  x"00",  x"29",  x"09",  x"7a",  x"87",  x"87", -- 00C8
         x"87",  x"53",  x"5f",  x"cb",  x"fa",  x"ed",  x"4b",  x"a2", -- 00D0
         x"b7",  x"cb",  x"49",  x"20",  x"16",  x"cd",  x"87",  x"f9", -- 00D8
         x"dd",  x"cb",  x"01",  x"5e",  x"20",  x"04",  x"cb",  x"71", -- 00E0
         x"20",  x"38",  x"78",  x"43",  x"cd",  x"68",  x"e1",  x"58", -- 00E8
         x"cd",  x"87",  x"f9",  x"cb",  x"41",  x"20",  x"12",  x"dd", -- 00F0
         x"cb",  x"01",  x"5e",  x"20",  x"04",  x"cb",  x"71",  x"20", -- 00F8
         x"2c",  x"cb",  x"51",  x"cc",  x"47",  x"e1",  x"c4",  x"5a", -- 0100
         x"e1",  x"cb",  x"69",  x"28",  x"8a",  x"f1",  x"dd",  x"77", -- 0108
         x"04",  x"d3",  x"86",  x"18",  x"82",  x"dd",  x"7e",  x"04", -- 0110
         x"f5",  x"dd",  x"cb",  x"04",  x"ff",  x"d3",  x"86",  x"c3", -- 0118
         x"b3",  x"d1",  x"78",  x"0f",  x"e5",  x"d5",  x"cd",  x"37", -- 0120
         x"e1",  x"d1",  x"e1",  x"18",  x"c3",  x"78",  x"e5",  x"d5", -- 0128
         x"cd",  x"37",  x"e1",  x"d1",  x"e1",  x"18",  x"d2",  x"e6", -- 0130
         x"09",  x"28",  x"2d",  x"ea",  x"66",  x"e1",  x"cb",  x"51", -- 0138
         x"28",  x"02",  x"ee",  x"09",  x"3d",  x"28",  x"13",  x"c5", -- 0140
         x"ed",  x"a0",  x"ed",  x"a0",  x"ed",  x"a0",  x"ed",  x"a0", -- 0148
         x"ed",  x"a0",  x"ed",  x"a0",  x"ed",  x"a0",  x"ed",  x"a0", -- 0150
         x"c1",  x"c9",  x"c5",  x"06",  x"08",  x"7e",  x"2f",  x"12", -- 0158
         x"23",  x"1c",  x"10",  x"f9",  x"c1",  x"c9",  x"3e",  x"ff", -- 0160
         x"12",  x"1c",  x"12",  x"1c",  x"12",  x"1c",  x"12",  x"1c", -- 0168
         x"12",  x"1c",  x"12",  x"1c",  x"12",  x"1c",  x"12",  x"c9", -- 0170
         x"ed",  x"5b",  x"a0",  x"b7",  x"21",  x"a2",  x"b7",  x"cb", -- 0178
         x"66",  x"28",  x"22",  x"cb",  x"a6",  x"fe",  x"30",  x"d8", -- 0180
         x"fe",  x"3a",  x"30",  x"04",  x"d6",  x"30",  x"18",  x"0a", -- 0188
         x"fe",  x"41",  x"d8",  x"cb",  x"af",  x"fe",  x"5b",  x"d0", -- 0190
         x"d6",  x"37",  x"21",  x"df",  x"b7",  x"be",  x"d0",  x"87", -- 0198
         x"2a",  x"dd",  x"b7",  x"18",  x"0c",  x"fe",  x"20",  x"30", -- 01A0
         x"18",  x"cb",  x"5e",  x"20",  x"14",  x"87",  x"2a",  x"b2", -- 01A8
         x"b7",  x"4f",  x"06",  x"00",  x"09",  x"7e",  x"23",  x"66", -- 01B0
         x"6f",  x"e9",  x"7b",  x"f6",  x"07",  x"3c",  x"5f",  x"18", -- 01B8
         x"09",  x"cd",  x"68",  x"e0",  x"d8",  x"77",  x"cd",  x"9c", -- 01C0
         x"e0",  x"1c",  x"3a",  x"9e",  x"b7",  x"3d",  x"bb",  x"d0", -- 01C8
         x"1e",  x"00",  x"14",  x"3a",  x"9f",  x"b7",  x"ba",  x"c0", -- 01D0
         x"2a",  x"a4",  x"b7",  x"e9",  x"2a",  x"99",  x"b7",  x"e9", -- 01D8
         x"7b",  x"a7",  x"28",  x"02",  x"1d",  x"c9",  x"7a",  x"a7", -- 01E0
         x"c8",  x"15",  x"3a",  x"9e",  x"b7",  x"3d",  x"5f",  x"c9", -- 01E8
         x"7a",  x"a7",  x"c8",  x"15",  x"c9",  x"21",  x"64",  x"e2", -- 01F0
         x"22",  x"a4",  x"b7",  x"c9",  x"21",  x"69",  x"e2",  x"18", -- 01F8
         x"f7",  x"cd",  x"e0",  x"e1",  x"d5",  x"cd",  x"68",  x"e0", -- 0200
         x"7e",  x"a7",  x"28",  x"29",  x"e5",  x"d5",  x"1c",  x"cd", -- 0208
         x"68",  x"e0",  x"30",  x"08",  x"1e",  x"00",  x"14",  x"cd", -- 0210
         x"68",  x"e0",  x"38",  x"10",  x"7e",  x"a7",  x"28",  x"0c", -- 0218
         x"42",  x"4b",  x"d1",  x"e3",  x"77",  x"cd",  x"9c",  x"e0", -- 0220
         x"50",  x"59",  x"18",  x"e1",  x"d1",  x"e1",  x"36",  x"00", -- 0228
         x"3e",  x"20",  x"cd",  x"9c",  x"e0",  x"d1",  x"c9",  x"d5", -- 0230
         x"3e",  x"20",  x"cd",  x"68",  x"e0",  x"46",  x"77",  x"cd", -- 0238
         x"9c",  x"e0",  x"78",  x"a7",  x"28",  x"0e",  x"1c",  x"cd", -- 0240
         x"68",  x"e0",  x"30",  x"f1",  x"1e",  x"00",  x"14",  x"cd", -- 0248
         x"68",  x"e0",  x"30",  x"e9",  x"d1",  x"c9",  x"3a",  x"9f", -- 0250
         x"b7",  x"16",  x"00",  x"f5",  x"cd",  x"78",  x"e2",  x"f1", -- 0258
         x"14",  x"3d",  x"20",  x"f7",  x"16",  x"00",  x"1e",  x"00", -- 0260
         x"c9",  x"dd",  x"7e",  x"04",  x"f5",  x"dd",  x"cb",  x"04", -- 0268
         x"ff",  x"d3",  x"86",  x"cd",  x"33",  x"d2",  x"18",  x"0d", -- 0270
         x"dd",  x"7e",  x"04",  x"f5",  x"dd",  x"cb",  x"04",  x"ff", -- 0278
         x"d3",  x"86",  x"cd",  x"7a",  x"d2",  x"f1",  x"dd",  x"77", -- 0280
         x"04",  x"d3",  x"86",  x"c9",  x"01",  x"0f",  x"0a",  x"21", -- 0288
         x"30",  x"00",  x"d5",  x"5c",  x"cd",  x"15",  x"f9",  x"3e", -- 0290
         x"1e",  x"cd",  x"a3",  x"e2",  x"3e",  x"03",  x"d3",  x"8c", -- 0298
         x"3e",  x"10",  x"d1",  x"47",  x"af",  x"cd",  x"ab",  x"e2", -- 02A0
         x"10",  x"fb",  x"c9",  x"3d",  x"c8",  x"f5",  x"f1",  x"18", -- 02A8
         x"fa",  x"01",  x"07",  x"03",  x"21",  x"24",  x"00",  x"d5", -- 02B0
         x"5c",  x"cd",  x"15",  x"f9",  x"d1",  x"c9",  x"21",  x"a3", -- 02B8
         x"b7",  x"7e",  x"e6",  x"07",  x"07",  x"07",  x"07",  x"4f", -- 02C0
         x"7e",  x"e6",  x"38",  x"0f",  x"0f",  x"0f",  x"b1",  x"4f", -- 02C8
         x"7e",  x"e6",  x"c0",  x"b1",  x"77",  x"c9",  x"7e",  x"c9", -- 02D0
         x"dd",  x"7e",  x"08",  x"ee",  x"20",  x"dd",  x"77",  x"08", -- 02D8
         x"c9",  x"fb",  x"f5",  x"3e",  x"23",  x"d3",  x"8f",  x"dd", -- 02E0
         x"36",  x"0d",  x"00",  x"18",  x"5a",  x"f5",  x"db",  x"8f", -- 02E8
         x"f5",  x"3e",  x"a7",  x"d3",  x"8f",  x"3e",  x"8f",  x"d3", -- 02F0
         x"8f",  x"f1",  x"fb",  x"fe",  x"14",  x"38",  x"48",  x"fe", -- 02F8
         x"78",  x"30",  x"44",  x"fe",  x"65",  x"30",  x"04",  x"c6", -- 0300
         x"be",  x"30",  x"06",  x"dd",  x"cb",  x"0c",  x"1e",  x"18", -- 0308
         x"36",  x"e5",  x"d5",  x"dd",  x"7e",  x"0c",  x"1f",  x"ee", -- 0310
         x"01",  x"dd",  x"6e",  x"0e",  x"dd",  x"66",  x"0f",  x"16", -- 0318
         x"00",  x"5f",  x"19",  x"7e",  x"dd",  x"cb",  x"08",  x"7e", -- 0320
         x"20",  x"07",  x"fe",  x"40",  x"fa",  x"31",  x"e3",  x"ee", -- 0328
         x"20",  x"57",  x"dd",  x"be",  x"0d",  x"20",  x"17",  x"21", -- 0330
         x"e0",  x"b7",  x"cd",  x"86",  x"e3",  x"dd",  x"be",  x"0a", -- 0338
         x"38",  x"1c",  x"dd",  x"34",  x"0a",  x"d1",  x"e1",  x"db", -- 0340
         x"89",  x"d3",  x"89",  x"f1",  x"ed",  x"4d",  x"dd",  x"36", -- 0348
         x"0a",  x"00",  x"fe",  x"16",  x"20",  x"09",  x"dd",  x"7e", -- 0350
         x"08",  x"ee",  x"80",  x"dd",  x"77",  x"08",  x"7a",  x"dd", -- 0358
         x"77",  x"0d",  x"dd",  x"cb",  x"08",  x"c6",  x"18",  x"dd", -- 0360
         x"b7",  x"dd",  x"cb",  x"08",  x"46",  x"c8",  x"dd",  x"7e", -- 0368
         x"0d",  x"37",  x"c9",  x"cd",  x"68",  x"e3",  x"d0",  x"dd", -- 0370
         x"cb",  x"08",  x"86",  x"c9",  x"cd",  x"68",  x"e3",  x"d0", -- 0378
         x"fe",  x"03",  x"37",  x"c8",  x"a7",  x"c9",  x"d5",  x"db", -- 0380
         x"88",  x"5f",  x"cb",  x"d7",  x"f3",  x"d3",  x"88",  x"56", -- 0388
         x"7b",  x"d3",  x"88",  x"fb",  x"7a",  x"d1",  x"c9",  x"f5", -- 0390
         x"e5",  x"d5",  x"c5",  x"21",  x"00",  x"a8",  x"cd",  x"86", -- 0398
         x"e3",  x"47",  x"0e",  x"80",  x"3e",  x"01",  x"ed",  x"79", -- 03A0
         x"db",  x"09",  x"5f",  x"a7",  x"28",  x"0e",  x"dd",  x"be", -- 03A8
         x"0d",  x"3e",  x"00",  x"20",  x"07",  x"21",  x"e0",  x"b7", -- 03B0
         x"cd",  x"86",  x"e3",  x"3c",  x"dd",  x"77",  x"0a",  x"7b", -- 03B8
         x"dd",  x"77",  x"0d",  x"a7",  x"28",  x"04",  x"dd",  x"cb", -- 03C0
         x"08",  x"c6",  x"26",  x"b8",  x"68",  x"cd",  x"86",  x"e3", -- 03C8
         x"ed",  x"79",  x"c1",  x"18",  x"48",  x"f5",  x"db",  x"90", -- 03D0
         x"fb",  x"2f",  x"e5",  x"d5",  x"e6",  x"3f",  x"28",  x"42", -- 03D8
         x"fe",  x"10",  x"38",  x"06",  x"e6",  x"30",  x"0f",  x"0f", -- 03E0
         x"ee",  x"0f",  x"c5",  x"4f",  x"06",  x"00",  x"db",  x"88", -- 03E8
         x"57",  x"f6",  x"04",  x"f3",  x"d3",  x"88",  x"2a",  x"f0", -- 03F0
         x"b7",  x"5e",  x"09",  x"6e",  x"3a",  x"e0",  x"b7",  x"67", -- 03F8
         x"7a",  x"d3",  x"88",  x"fb",  x"c1",  x"3e",  x"4f",  x"d3", -- 0400
         x"92",  x"7d",  x"a7",  x"28",  x"10",  x"dd",  x"be",  x"0d", -- 0408
         x"28",  x"28",  x"dd",  x"77",  x"0d",  x"af",  x"dd",  x"cb", -- 0410
         x"08",  x"c6",  x"dd",  x"77",  x"0a",  x"d1",  x"e1",  x"f1", -- 0418
         x"ed",  x"4d",  x"dd",  x"be",  x"0a",  x"3c",  x"30",  x"f2", -- 0420
         x"21",  x"9e",  x"ed",  x"f3",  x"cd",  x"4f",  x"f5",  x"fb", -- 0428
         x"af",  x"dd",  x"77",  x"0d",  x"dd",  x"cb",  x"08",  x"86", -- 0430
         x"18",  x"e0",  x"7c",  x"87",  x"87",  x"bb",  x"30",  x"01", -- 0438
         x"7b",  x"67",  x"dd",  x"7e",  x"0a",  x"bc",  x"3c",  x"38", -- 0440
         x"d1",  x"7c",  x"93",  x"18",  x"c9",  x"dd",  x"36",  x"03", -- 0448
         x"01",  x"f3",  x"db",  x"88",  x"f6",  x"40",  x"e6",  x"df", -- 0450
         x"d3",  x"88",  x"fb",  x"2a",  x"a4",  x"b7",  x"22",  x"cf", -- 0458
         x"b7",  x"cd",  x"8c",  x"f3",  x"22",  x"cd",  x"b7",  x"cd", -- 0460
         x"f5",  x"e1",  x"3e",  x"03",  x"d3",  x"8c",  x"d3",  x"8d", -- 0468
         x"dd",  x"cb",  x"08",  x"8e",  x"18",  x"1d",  x"dd",  x"36", -- 0470
         x"02",  x"fe",  x"cd",  x"0f",  x"d0",  x"2a",  x"cd",  x"b7", -- 0478
         x"22",  x"b9",  x"b7",  x"2a",  x"cf",  x"b7",  x"22",  x"a4", -- 0480
         x"b7",  x"db",  x"88",  x"e6",  x"9f",  x"d3",  x"88",  x"dd", -- 0488
         x"cb",  x"08",  x"86",  x"dd",  x"cb",  x"01",  x"5e",  x"28", -- 0490
         x"06",  x"db",  x"89",  x"cb",  x"ff",  x"d3",  x"89",  x"dd", -- 0498
         x"cb",  x"08",  x"4e",  x"20",  x"fa",  x"db",  x"88",  x"6f", -- 04A0
         x"cb",  x"d7",  x"f3",  x"d3",  x"88",  x"3a",  x"db",  x"b7", -- 04A8
         x"e6",  x"60",  x"f6",  x"07",  x"d3",  x"8e",  x"3a",  x"dc", -- 04B0
         x"b7",  x"d3",  x"8e",  x"7d",  x"d3",  x"88",  x"fb",  x"c9", -- 04B8
         x"11",  x"80",  x"b7",  x"af",  x"1d",  x"12",  x"20",  x"fc", -- 04C0
         x"c9",  x"e5",  x"21",  x"3a",  x"e5",  x"e3",  x"e5",  x"f3", -- 04C8
         x"e1",  x"e1",  x"e1",  x"23",  x"e5",  x"2b",  x"3b",  x"3b", -- 04D0
         x"3b",  x"3b",  x"fb",  x"f5",  x"7e",  x"fe",  x"0c",  x"38", -- 04D8
         x"03",  x"f1",  x"e1",  x"c9",  x"87",  x"c6",  x"08",  x"6f", -- 04E0
         x"cd",  x"90",  x"ed",  x"b5",  x"6f",  x"26",  x"a9",  x"7e", -- 04E8
         x"23",  x"66",  x"6f",  x"f1",  x"e3",  x"e5",  x"d5",  x"c5", -- 04F0
         x"f5",  x"26",  x"a9",  x"cd",  x"90",  x"ed",  x"f6",  x"01", -- 04F8
         x"6f",  x"5e",  x"16",  x"b8",  x"1a",  x"2c",  x"77",  x"2c", -- 0500
         x"7e",  x"12",  x"57",  x"7b",  x"1e",  x"00",  x"fe",  x"05", -- 0508
         x"20",  x"02",  x"1e",  x"80",  x"fe",  x"07",  x"38",  x"05", -- 0510
         x"0e",  x"80",  x"47",  x"ed",  x"51",  x"db",  x"88",  x"e6", -- 0518
         x"7f",  x"d3",  x"88",  x"21",  x"05",  x"b8",  x"dd",  x"7e", -- 0520
         x"04",  x"e6",  x"80",  x"b6",  x"77",  x"dd",  x"7e",  x"04", -- 0528
         x"e6",  x"7f",  x"b3",  x"dd",  x"77",  x"04",  x"d3",  x"86", -- 0530
         x"18",  x"39",  x"e5",  x"d5",  x"c5",  x"f5",  x"21",  x"02", -- 0538
         x"b8",  x"56",  x"cd",  x"02",  x"f1",  x"26",  x"a9",  x"cd", -- 0540
         x"90",  x"ed",  x"f6",  x"02",  x"6f",  x"56",  x"2d",  x"7e", -- 0548
         x"6f",  x"fe",  x"05",  x"28",  x"09",  x"cd",  x"02",  x"f1", -- 0550
         x"3a",  x"05",  x"b8",  x"e6",  x"01",  x"57",  x"21",  x"05", -- 0558
         x"b8",  x"7e",  x"72",  x"e6",  x"80",  x"dd",  x"7e",  x"04", -- 0560
         x"cb",  x"bf",  x"28",  x"02",  x"cb",  x"ff",  x"dd",  x"77", -- 0568
         x"04",  x"d3",  x"86",  x"c3",  x"97",  x"e0",  x"cd",  x"c9", -- 0570
         x"e4",  x"00",  x"c9",  x"cd",  x"c9",  x"e4",  x"01",  x"c9", -- 0578
         x"cd",  x"c9",  x"e4",  x"02",  x"c9",  x"cd",  x"c9",  x"e4", -- 0580
         x"03",  x"c9",  x"cd",  x"c9",  x"e4",  x"04",  x"c9",  x"cd", -- 0588
         x"c9",  x"e4",  x"05",  x"c9",  x"f5",  x"3e",  x"87",  x"d3", -- 0590
         x"8d",  x"dd",  x"7e",  x"00",  x"d3",  x"8d",  x"dd",  x"36", -- 0598
         x"00",  x"00",  x"18",  x"0e",  x"f5",  x"db",  x"8e",  x"dd", -- 05A0
         x"77",  x"00",  x"3e",  x"07",  x"d3",  x"8e",  x"3e",  x"a3", -- 05A8
         x"d3",  x"8e",  x"f1",  x"fb",  x"ed",  x"4d",  x"78",  x"d6", -- 05B0
         x"09",  x"38",  x"48",  x"fe",  x"1f",  x"30",  x"44",  x"07", -- 05B8
         x"4f",  x"06",  x"00",  x"eb",  x"21",  x"91",  x"fd",  x"c3", -- 05C0
         x"b7",  x"c8",  x"e5",  x"21",  x"a3",  x"b7",  x"cd",  x"1d", -- 05C8
         x"eb",  x"e1",  x"c9",  x"7e",  x"fe",  x"df",  x"d8",  x"fe", -- 05D0
         x"e3",  x"d0",  x"fe",  x"e1",  x"ca",  x"45",  x"e9",  x"3a", -- 05D8
         x"fd",  x"03",  x"a7",  x"20",  x"1e",  x"3c",  x"32",  x"fd", -- 05E0
         x"03",  x"cd",  x"ca",  x"e5",  x"32",  x"7e",  x"03",  x"7e", -- 05E8
         x"fe",  x"df",  x"28",  x"1a",  x"fe",  x"e2",  x"28",  x"0e", -- 05F0
         x"cd",  x"bd",  x"c8",  x"cd",  x"1c",  x"ea",  x"7e",  x"fe", -- 05F8
         x"3b",  x"28",  x"3b",  x"c3",  x"48",  x"c3",  x"cd",  x"bd", -- 0600
         x"c8",  x"cd",  x"0d",  x"ea",  x"18",  x"f0",  x"cd",  x"bd", -- 0608
         x"c8",  x"cd",  x"fb",  x"e9",  x"7e",  x"fe",  x"3b",  x"28", -- 0610
         x"25",  x"cd",  x"cc",  x"c8",  x"2c",  x"fe",  x"e0",  x"20", -- 0618
         x"e2",  x"cd",  x"bd",  x"c8",  x"cd",  x"1c",  x"ea",  x"cd", -- 0620
         x"cc",  x"c8",  x"3b",  x"cd",  x"03",  x"cb",  x"3a",  x"7e", -- 0628
         x"03",  x"e5",  x"21",  x"a3",  x"b7",  x"cd",  x"22",  x"eb", -- 0630
         x"e1",  x"c1",  x"c9",  x"c5",  x"18",  x"ab",  x"cd",  x"bd", -- 0638
         x"c8",  x"18",  x"e8",  x"cd",  x"cc",  x"c8",  x"28",  x"cd", -- 0640
         x"21",  x"d4",  x"f5",  x"cd",  x"d6",  x"c8",  x"cd",  x"3a", -- 0648
         x"cd",  x"cd",  x"db",  x"c8",  x"f1",  x"e5",  x"f5",  x"cd", -- 0650
         x"30",  x"d3",  x"23",  x"23",  x"5e",  x"23",  x"56",  x"c1", -- 0658
         x"c5",  x"f5",  x"d5",  x"4f",  x"af",  x"b9",  x"28",  x"0c", -- 0660
         x"b8",  x"28",  x"09",  x"79",  x"05",  x"28",  x"05",  x"81", -- 0668
         x"38",  x"2b",  x"10",  x"fb",  x"47",  x"0e",  x"00",  x"c5", -- 0670
         x"cd",  x"e1",  x"d1",  x"c1",  x"c1",  x"c5",  x"cd",  x"7e", -- 0678
         x"d1",  x"e1",  x"e3",  x"7c",  x"e1",  x"e3",  x"6f",  x"24", -- 0680
         x"25",  x"e5",  x"c5",  x"28",  x"07",  x"cd",  x"f2",  x"d2", -- 0688
         x"c1",  x"e1",  x"18",  x"f4",  x"c1",  x"e1",  x"d1",  x"cd", -- 0690
         x"02",  x"d3",  x"c3",  x"a9",  x"d1",  x"1e",  x"1c",  x"c3", -- 0698
         x"56",  x"c3",  x"e5",  x"21",  x"0a",  x"00",  x"22",  x"54", -- 06A0
         x"03",  x"2a",  x"5f",  x"03",  x"f5",  x"e5",  x"23",  x"23", -- 06A8
         x"7e",  x"23",  x"66",  x"6f",  x"22",  x"4e",  x"03",  x"22", -- 06B0
         x"52",  x"03",  x"ed",  x"5b",  x"d7",  x"03",  x"1b",  x"1b", -- 06B8
         x"e1",  x"e5",  x"7e",  x"23",  x"66",  x"6f",  x"cd",  x"89", -- 06C0
         x"c6",  x"e3",  x"20",  x"f4",  x"d1",  x"23",  x"23",  x"7e", -- 06C8
         x"23",  x"66",  x"6f",  x"22",  x"50",  x"03",  x"06",  x"04", -- 06D0
         x"f1",  x"21",  x"4e",  x"03",  x"e3",  x"28",  x"20",  x"cd", -- 06D8
         x"86",  x"c9",  x"f5",  x"7a",  x"b3",  x"ca",  x"67",  x"c9", -- 06E0
         x"f1",  x"e3",  x"73",  x"23",  x"72",  x"23",  x"28",  x"0f", -- 06E8
         x"f5",  x"05",  x"28",  x"07",  x"f1",  x"e3",  x"cd",  x"d6", -- 06F0
         x"c8",  x"18",  x"e2",  x"f1",  x"c2",  x"48",  x"c3",  x"2a", -- 06F8
         x"50",  x"03",  x"ed",  x"5b",  x"4e",  x"03",  x"cd",  x"89", -- 0700
         x"c6",  x"da",  x"67",  x"c9",  x"2a",  x"5f",  x"03",  x"cd", -- 0708
         x"be",  x"c4",  x"38",  x"04",  x"28",  x"cf",  x"18",  x"f7", -- 0710
         x"e1",  x"c5",  x"ed",  x"5b",  x"50",  x"03",  x"21",  x"00", -- 0718
         x"00",  x"22",  x"50",  x"03",  x"60",  x"69",  x"4e",  x"23", -- 0720
         x"46",  x"78",  x"b1",  x"28",  x"b8",  x"23",  x"7e",  x"23", -- 0728
         x"66",  x"6f",  x"cd",  x"89",  x"c6",  x"2a",  x"50",  x"03", -- 0730
         x"23",  x"22",  x"50",  x"03",  x"20",  x"e6",  x"23",  x"23", -- 0738
         x"29",  x"23",  x"ed",  x"5b",  x"d7",  x"03",  x"19",  x"38", -- 0740
         x"c0",  x"cd",  x"27",  x"c3",  x"22",  x"d7",  x"03",  x"af", -- 0748
         x"2b",  x"77",  x"2b",  x"77",  x"1b",  x"1b",  x"eb",  x"73", -- 0750
         x"23",  x"72",  x"23",  x"3d",  x"77",  x"23",  x"77",  x"23", -- 0758
         x"eb",  x"2a",  x"52",  x"03",  x"22",  x"4e",  x"03",  x"e1", -- 0760
         x"4e",  x"23",  x"46",  x"23",  x"c5",  x"01",  x"4e",  x"03", -- 0768
         x"7e",  x"12",  x"0a",  x"77",  x"23",  x"13",  x"03",  x"7e", -- 0770
         x"12",  x"0a",  x"77",  x"13",  x"2a",  x"4e",  x"03",  x"ed", -- 0778
         x"4b",  x"54",  x"03",  x"09",  x"22",  x"4e",  x"03",  x"2a", -- 0780
         x"50",  x"03",  x"2b",  x"7c",  x"b5",  x"22",  x"50",  x"03", -- 0788
         x"20",  x"d5",  x"12",  x"e1",  x"2a",  x"5f",  x"03",  x"e5", -- 0790
         x"e1",  x"4e",  x"23",  x"46",  x"23",  x"c5",  x"7e",  x"23", -- 0798
         x"a6",  x"3c",  x"28",  x"26",  x"23",  x"7e",  x"b7",  x"28", -- 07A0
         x"ef",  x"fe",  x"88",  x"28",  x"2a",  x"fe",  x"8c",  x"28", -- 07A8
         x"26",  x"fe",  x"8b",  x"28",  x"08",  x"fe",  x"d4",  x"28", -- 07B0
         x"04",  x"fe",  x"a9",  x"20",  x"e7",  x"cd",  x"87",  x"c9", -- 07B8
         x"7b",  x"b2",  x"c4",  x"eb",  x"e7",  x"c4",  x"1c",  x"e8", -- 07C0
         x"18",  x"db",  x"2b",  x"22",  x"d7",  x"03",  x"2b",  x"77", -- 07C8
         x"2b",  x"77",  x"e1",  x"e1",  x"c3",  x"8a",  x"c4",  x"cd", -- 07D0
         x"87",  x"c9",  x"7b",  x"b2",  x"28",  x"c7",  x"cd",  x"eb", -- 07D8
         x"e7",  x"c4",  x"1c",  x"e8",  x"7e",  x"fe",  x"2c",  x"20", -- 07E0
         x"bc",  x"18",  x"ec",  x"e5",  x"d5",  x"11",  x"ff",  x"ff", -- 07E8
         x"cd",  x"bb",  x"c4",  x"d1",  x"03",  x"03",  x"03",  x"03", -- 07F0
         x"60",  x"69",  x"ed",  x"4b",  x"52",  x"03",  x"7e",  x"23", -- 07F8
         x"e5",  x"b6",  x"28",  x"15",  x"7e",  x"2b",  x"6e",  x"67", -- 0800
         x"cd",  x"89",  x"c6",  x"28",  x"0a",  x"2a",  x"54",  x"03", -- 0808
         x"09",  x"44",  x"4d",  x"e1",  x"23",  x"18",  x"e7",  x"af", -- 0810
         x"3d",  x"e1",  x"e1",  x"c9",  x"c5",  x"eb",  x"2a",  x"d7", -- 0818
         x"03",  x"ed",  x"52",  x"e5",  x"c1",  x"62",  x"6b",  x"1b", -- 0820
         x"1a",  x"fe",  x"2c",  x"28",  x"0b",  x"fe",  x"3a",  x"30", -- 0828
         x"07",  x"c5",  x"d5",  x"ed",  x"b0",  x"d1",  x"18",  x"ec", -- 0830
         x"eb",  x"d1",  x"e5",  x"c5",  x"af",  x"06",  x"98",  x"cd", -- 0838
         x"ae",  x"d6",  x"cd",  x"34",  x"d8",  x"c1",  x"d1",  x"23", -- 0840
         x"13",  x"7e",  x"b7",  x"28",  x"0f",  x"c5",  x"e5",  x"eb", -- 0848
         x"09",  x"54",  x"5d",  x"2b",  x"ed",  x"b8",  x"e1",  x"ed", -- 0850
         x"a0",  x"c1",  x"18",  x"ed",  x"d5",  x"ed",  x"5b",  x"5f", -- 0858
         x"03",  x"cd",  x"93",  x"c4",  x"23",  x"7e",  x"23",  x"b6", -- 0860
         x"20",  x"fa",  x"eb",  x"73",  x"23",  x"72",  x"13",  x"13", -- 0868
         x"ed",  x"53",  x"d7",  x"03",  x"e1",  x"54",  x"5d",  x"7e", -- 0870
         x"b7",  x"23",  x"20",  x"fb",  x"c1",  x"e3",  x"c5",  x"eb", -- 0878
         x"c9",  x"c8",  x"cd",  x"86",  x"c9",  x"ca",  x"42",  x"c4", -- 0880
         x"cd",  x"d6",  x"c8",  x"d5",  x"cd",  x"86",  x"c9",  x"e1", -- 0888
         x"c0",  x"eb",  x"e5",  x"cd",  x"bb",  x"c4",  x"30",  x"0a", -- 0890
         x"d1",  x"f5",  x"c5",  x"cd",  x"be",  x"c4",  x"c1",  x"da", -- 0898
         x"50",  x"c4",  x"c3",  x"4d",  x"c4",  x"cd",  x"be",  x"c8", -- 08A0
         x"20",  x"0f",  x"cd",  x"68",  x"e3",  x"30",  x"fb",  x"fe", -- 08A8
         x"03",  x"c8",  x"fe",  x"0a",  x"20",  x"f4",  x"c3",  x"e4", -- 08B0
         x"dd",  x"cd",  x"21",  x"d4",  x"4f",  x"3e",  x"10",  x"cd", -- 08B8
         x"a3",  x"e2",  x"cd",  x"68",  x"e3",  x"30",  x"0a",  x"fe", -- 08C0
         x"03",  x"c8",  x"fe",  x"0a",  x"20",  x"03",  x"c3",  x"e4", -- 08C8
         x"dd",  x"0d",  x"20",  x"e9",  x"c9",  x"06",  x"01",  x"cd", -- 08D0
         x"be",  x"c8",  x"28",  x"04",  x"cd",  x"21",  x"d4",  x"47", -- 08D8
         x"3e",  x"07",  x"1e",  x"00",  x"cd",  x"2d",  x"f0",  x"10", -- 08E0
         x"f7",  x"c9",  x"cd",  x"d6",  x"c8",  x"c3",  x"21",  x"d4", -- 08E8
         x"cd",  x"be",  x"c8",  x"28",  x"31",  x"cd",  x"21",  x"d4", -- 08F0
         x"47",  x"c5",  x"cd",  x"ea",  x"e8",  x"57",  x"d5",  x"cd", -- 08F8
         x"ea",  x"e8",  x"d1",  x"5f",  x"d5",  x"cd",  x"ea",  x"e8", -- 0900
         x"d1",  x"e3",  x"6b",  x"93",  x"38",  x"34",  x"3c",  x"5f", -- 0908
         x"7a",  x"94",  x"38",  x"2e",  x"3c",  x"57",  x"cd",  x"83", -- 0910
         x"f0",  x"3a",  x"9b",  x"b7",  x"cd",  x"f7",  x"f7",  x"cd", -- 0918
         x"a0",  x"f0",  x"38",  x"1e",  x"e1",  x"c9",  x"e5",  x"21", -- 0920
         x"00",  x"01",  x"11",  x"28",  x"1e",  x"18",  x"e7",  x"cd", -- 0928
         x"6c",  x"c9",  x"d5",  x"cd",  x"ea",  x"e8",  x"e3",  x"11", -- 0930
         x"00",  x"80",  x"19",  x"38",  x"05",  x"cb",  x"74",  x"ca", -- 0938
         x"d8",  x"e9",  x"c3",  x"48",  x"c3",  x"3a",  x"fd",  x"03", -- 0940
         x"cb",  x"4f",  x"cb",  x"cf",  x"32",  x"fd",  x"03",  x"20", -- 0948
         x"f1",  x"d5",  x"e5",  x"cd",  x"83",  x"f0",  x"21",  x"9c", -- 0950
         x"b7",  x"22",  x"f6",  x"b9",  x"11",  x"ec",  x"b9",  x"01", -- 0958
         x"06",  x"00",  x"ed",  x"b0",  x"21",  x"00",  x"00",  x"22", -- 0960
         x"9c",  x"b7",  x"21",  x"28",  x"20",  x"22",  x"9e",  x"b7", -- 0968
         x"cd",  x"a0",  x"f0",  x"e1",  x"cd",  x"a5",  x"e9",  x"cd", -- 0970
         x"db",  x"c8",  x"cd",  x"cc",  x"c8",  x"3b",  x"7e",  x"fe", -- 0978
         x"df",  x"38",  x"1d",  x"fe",  x"e3",  x"30",  x"19",  x"cd", -- 0980
         x"3b",  x"e6",  x"e5",  x"cd",  x"83",  x"f0",  x"21",  x"ec", -- 0988
         x"b9",  x"11",  x"9c",  x"b7",  x"01",  x"06",  x"00",  x"ed", -- 0990
         x"b0",  x"cd",  x"a0",  x"f0",  x"e1",  x"d1",  x"c1",  x"c9", -- 0998
         x"cd",  x"03",  x"cb",  x"18",  x"e5",  x"cd",  x"bd",  x"c8", -- 09A0
         x"cd",  x"cc",  x"c8",  x"28",  x"cd",  x"21",  x"d4",  x"57", -- 09A8
         x"e5",  x"21",  x"9f",  x"b7",  x"cd",  x"1d",  x"eb",  x"e1", -- 09B0
         x"3d",  x"ba",  x"38",  x"3c",  x"d5",  x"cd",  x"ea",  x"e8", -- 09B8
         x"d1",  x"4f",  x"e5",  x"21",  x"9e",  x"b7",  x"cd",  x"1d", -- 09C0
         x"eb",  x"e1",  x"3d",  x"b9",  x"38",  x"2a",  x"79",  x"e5", -- 09C8
         x"21",  x"a0",  x"b7",  x"cd",  x"22",  x"eb",  x"7a",  x"23", -- 09D0
         x"cd",  x"22",  x"eb",  x"e1",  x"c9",  x"e5",  x"cd",  x"68", -- 09D8
         x"e3",  x"30",  x"0f",  x"3e",  x"01",  x"cd",  x"7b",  x"d1", -- 09E0
         x"cd",  x"e4",  x"dd",  x"2a",  x"c2",  x"03",  x"77",  x"c3", -- 09E8
         x"a9",  x"d1",  x"af",  x"cd",  x"7b",  x"d1",  x"18",  x"f7", -- 09F0
         x"c3",  x"48",  x"c3",  x"cd",  x"21",  x"d4",  x"fe",  x"20", -- 09F8
         x"30",  x"66",  x"87",  x"87",  x"87",  x"57",  x"cd",  x"ca", -- 0A00
         x"e5",  x"e6",  x"07",  x"18",  x"1c",  x"cd",  x"be",  x"c8", -- 0A08
         x"28",  x"56",  x"cd",  x"fb",  x"e9",  x"cd",  x"be",  x"c8", -- 0A10
         x"c8",  x"cd",  x"d6",  x"c8",  x"cd",  x"21",  x"d4",  x"fe", -- 0A18
         x"08",  x"30",  x"45",  x"57",  x"cd",  x"ca",  x"e5",  x"e6", -- 0A20
         x"f8",  x"b2",  x"e5",  x"21",  x"a3",  x"b7",  x"18",  x"a8", -- 0A28
         x"1e",  x"2f",  x"01",  x"1e",  x"30",  x"d5",  x"cd",  x"6c", -- 0A30
         x"c9",  x"e5",  x"7b",  x"21",  x"d3",  x"b7",  x"cd",  x"22", -- 0A38
         x"eb",  x"7a",  x"23",  x"cd",  x"22",  x"eb",  x"e3",  x"cd", -- 0A40
         x"ea",  x"e8",  x"e3",  x"23",  x"cd",  x"22",  x"eb",  x"e1", -- 0A48
         x"cd",  x"be",  x"c8",  x"28",  x"0e",  x"cd",  x"ea",  x"e8", -- 0A50
         x"17",  x"17",  x"17",  x"e5",  x"21",  x"d6",  x"b7",  x"cd", -- 0A58
         x"22",  x"eb",  x"e1",  x"d1",  x"cd",  x"2d",  x"f0",  x"d0", -- 0A60
         x"c3",  x"67",  x"c9",  x"cd",  x"21",  x"d4",  x"e5",  x"21", -- 0A68
         x"82",  x"b7",  x"06",  x"04",  x"cd",  x"22",  x"eb",  x"23", -- 0A70
         x"e3",  x"05",  x"28",  x"08",  x"c5",  x"cd",  x"ea",  x"e8", -- 0A78
         x"c1",  x"e3",  x"18",  x"f0",  x"cd",  x"be",  x"c8",  x"28", -- 0A80
         x"16",  x"cd",  x"ea",  x"e8",  x"e3",  x"cd",  x"22",  x"eb", -- 0A88
         x"23",  x"e3",  x"cd",  x"be",  x"c8",  x"28",  x"08",  x"cd", -- 0A90
         x"ea",  x"e8",  x"e3",  x"cd",  x"22",  x"eb",  x"e3",  x"1e", -- 0A98
         x"35",  x"c1",  x"c3",  x"2d",  x"f0",  x"cd",  x"36",  x"cd", -- 0AA0
         x"cd",  x"d6",  x"c8",  x"e5",  x"cd",  x"30",  x"d3",  x"28", -- 0AA8
         x"b7",  x"47",  x"23",  x"23",  x"5e",  x"23",  x"56",  x"e1", -- 0AB0
         x"d5",  x"c5",  x"cd",  x"3a",  x"cd",  x"cd",  x"db",  x"c8", -- 0AB8
         x"c1",  x"d1",  x"e5",  x"d5",  x"c5",  x"cd",  x"30",  x"d3", -- 0AC0
         x"28",  x"9e",  x"23",  x"23",  x"4e",  x"23",  x"66",  x"69", -- 0AC8
         x"c1",  x"4f",  x"d1",  x"e5",  x"c5",  x"d5",  x"1a",  x"be", -- 0AD0
         x"28",  x"0f",  x"23",  x"0d",  x"20",  x"f9",  x"af",  x"e1", -- 0AD8
         x"e1",  x"e1",  x"11",  x"f3",  x"cd",  x"d5",  x"c3",  x"c0", -- 0AE0
         x"d0",  x"23",  x"e5",  x"2b",  x"23",  x"0d",  x"28",  x"0e", -- 0AE8
         x"13",  x"05",  x"28",  x"11",  x"1a",  x"be",  x"28",  x"f4", -- 0AF0
         x"e1",  x"d1",  x"c1",  x"0d",  x"18",  x"d6",  x"13",  x"05", -- 0AF8
         x"e1",  x"20",  x"db",  x"18",  x"01",  x"e1",  x"d1",  x"d1", -- 0B00
         x"d1",  x"a7",  x"ed",  x"52",  x"7d",  x"18",  x"d3",  x"cd", -- 0B08
         x"21",  x"d4",  x"fe",  x"10",  x"d2",  x"b7",  x"eb",  x"1e", -- 0B10
         x"39",  x"01",  x"1e",  x"3a",  x"01",  x"1e",  x"29",  x"c3", -- 0B18
         x"2d",  x"f0",  x"1e",  x"28",  x"18",  x"f9",  x"cd",  x"21", -- 0B20
         x"d4",  x"f5",  x"cd",  x"ea",  x"e8",  x"57",  x"f1",  x"e5", -- 0B28
         x"6f",  x"3e",  x"02",  x"1e",  x"26",  x"cd",  x"2d",  x"f0", -- 0B30
         x"e1",  x"c9",  x"cd",  x"36",  x"cd",  x"cd",  x"6f",  x"c9", -- 0B38
         x"e5",  x"7b",  x"21",  x"d3",  x"b7",  x"cd",  x"22",  x"eb", -- 0B40
         x"7a",  x"23",  x"cd",  x"22",  x"eb",  x"23",  x"e3",  x"0e", -- 0B48
         x"00",  x"7e",  x"fe",  x"2c",  x"20",  x"0a",  x"cd",  x"ea", -- 0B50
         x"e8",  x"e3",  x"cd",  x"22",  x"eb",  x"e3",  x"0e",  x"ff", -- 0B58
         x"cd",  x"db",  x"c8",  x"d1",  x"e3",  x"11",  x"f3",  x"cd", -- 0B60
         x"d5",  x"e5",  x"1e",  x"2f",  x"cd",  x"2d",  x"f0",  x"da", -- 0B68
         x"67",  x"c9",  x"f5",  x"dd",  x"cb",  x"01",  x"5e",  x"28", -- 0B70
         x"20",  x"f1",  x"06",  x"00",  x"28",  x"19",  x"21",  x"d6", -- 0B78
         x"b7",  x"cd",  x"22",  x"eb",  x"0f",  x"0f",  x"0f",  x"e6", -- 0B80
         x"0f",  x"20",  x"02",  x"3e",  x"08",  x"47",  x"1e",  x"30", -- 0B88
         x"cd",  x"2d",  x"f0",  x"0c",  x"28",  x"01",  x"41",  x"78", -- 0B90
         x"06",  x"f1",  x"18",  x"65",  x"cd",  x"e1",  x"cd",  x"e3", -- 0B98
         x"11",  x"f3",  x"cd",  x"d5",  x"cd",  x"6f",  x"c9",  x"e5", -- 0BA0
         x"21",  x"00",  x"80",  x"19",  x"38",  x"09",  x"cb",  x"74", -- 0BA8
         x"20",  x"05",  x"cd",  x"1d",  x"eb",  x"18",  x"4a",  x"c3", -- 0BB0
         x"48",  x"c3",  x"79",  x"fe",  x"62",  x"28",  x"dd",  x"fe", -- 0BB8
         x"6e",  x"ca",  x"3a",  x"eb",  x"fe",  x"7c",  x"28",  x"1a", -- 0BC0
         x"fe",  x"76",  x"28",  x"39",  x"d6",  x"3e",  x"38",  x"e7", -- 0BC8
         x"fe",  x"07",  x"30",  x"e3",  x"eb",  x"01",  x"89",  x"fd", -- 0BD0
         x"e1",  x"6f",  x"09",  x"4e",  x"23",  x"66",  x"69",  x"e5", -- 0BD8
         x"eb",  x"c9",  x"cd",  x"e1",  x"cd",  x"e3",  x"11",  x"f3", -- 0BE0
         x"cd",  x"d5",  x"cd",  x"24",  x"d4",  x"e5",  x"a7",  x"3e", -- 0BE8
         x"00",  x"20",  x"06",  x"21",  x"9d",  x"b7",  x"cd",  x"1d", -- 0BF0
         x"eb",  x"47",  x"21",  x"a1",  x"b7",  x"cd",  x"1d",  x"eb", -- 0BF8
         x"80",  x"e1",  x"c3",  x"c0",  x"d0",  x"e3",  x"3e",  x"01", -- 0C00
         x"cd",  x"7b",  x"d1",  x"cd",  x"83",  x"f0",  x"ed",  x"5b", -- 0C08
         x"a0",  x"b7",  x"cd",  x"68",  x"e0",  x"7e",  x"cd",  x"a0", -- 0C10
         x"f0",  x"c3",  x"eb",  x"e9",  x"0e",  x"00",  x"7e",  x"fe", -- 0C18
         x"49",  x"28",  x"05",  x"0c",  x"fe",  x"4f",  x"20",  x"8f", -- 0C20
         x"c5",  x"23",  x"7e",  x"fe",  x"23",  x"20",  x"88",  x"23", -- 0C28
         x"cd",  x"21",  x"d4",  x"e6",  x"03",  x"c1",  x"c8",  x"e5", -- 0C30
         x"17",  x"81",  x"f5",  x"3d",  x"47",  x"3e",  x"ff",  x"17", -- 0C38
         x"10",  x"fd",  x"21",  x"07",  x"03",  x"a6",  x"77",  x"f1", -- 0C40
         x"e1",  x"cb",  x"f7",  x"d5",  x"5f",  x"16",  x"03",  x"cd", -- 0C48
         x"0e",  x"e0",  x"d1",  x"c9",  x"cd",  x"e1",  x"cd",  x"e5", -- 0C50
         x"11",  x"f3",  x"cd",  x"d5",  x"cd",  x"6f",  x"c9",  x"7b", -- 0C58
         x"3d",  x"b2",  x"3e",  x"00",  x"20",  x"9c",  x"db",  x"90", -- 0C60
         x"2f",  x"57",  x"e6",  x"0f",  x"1f",  x"30",  x"02",  x"f6", -- 0C68
         x"10",  x"1f",  x"30",  x"02",  x"f6",  x"04",  x"5f",  x"3e", -- 0C70
         x"30",  x"a2",  x"b3",  x"18",  x"85",  x"ed",  x"5f",  x"32", -- 0C78
         x"1d",  x"03",  x"c9",  x"7e",  x"23",  x"fe",  x"49",  x"28", -- 0C80
         x"19",  x"fe",  x"4f",  x"20",  x"a0",  x"cd",  x"25",  x"de", -- 0C88
         x"cd",  x"c8",  x"dd",  x"c8",  x"3e",  x"d5",  x"cd",  x"b2", -- 0C90
         x"dc",  x"21",  x"ea",  x"03",  x"af",  x"cd",  x"d5",  x"dd", -- 0C98
         x"e1",  x"c9",  x"cd",  x"5f",  x"de",  x"3a",  x"09",  x"03", -- 0CA0
         x"e6",  x"03",  x"c8",  x"3e",  x"d5",  x"cd",  x"b2",  x"dc", -- 0CA8
         x"21",  x"ea",  x"03",  x"cd",  x"e4",  x"dd",  x"e1",  x"c9", -- 0CB0
         x"01",  x"3e",  x"04",  x"18",  x"03",  x"01",  x"3f",  x"03", -- 0CB8
         x"c5",  x"cd",  x"6c",  x"c9",  x"c1",  x"c5",  x"e5",  x"21", -- 0CC0
         x"82",  x"b7",  x"7b",  x"cd",  x"22",  x"eb",  x"23",  x"7a", -- 0CC8
         x"cd",  x"22",  x"eb",  x"23",  x"05",  x"ca",  x"4f",  x"ea", -- 0CD0
         x"e3",  x"c5",  x"cd",  x"d6",  x"c8",  x"cd",  x"6c",  x"c9", -- 0CD8
         x"c1",  x"e3",  x"18",  x"e6",  x"cd",  x"be",  x"c8",  x"3e", -- 0CE0
         x"ff",  x"c4",  x"21",  x"d4",  x"e5",  x"cd",  x"83",  x"f0", -- 0CE8
         x"cd",  x"d7",  x"fb",  x"da",  x"83",  x"f8",  x"3e",  x"fe", -- 0CF0
         x"cd",  x"d7",  x"fb",  x"cd",  x"db",  x"f4",  x"cd",  x"a0", -- 0CF8
         x"f0",  x"e1",  x"c9",  x"cd",  x"be",  x"c8",  x"28",  x"16", -- 0D00
         x"cd",  x"3a",  x"cd",  x"e5",  x"3e",  x"0c",  x"cd",  x"56", -- 0D08
         x"ed",  x"eb",  x"cd",  x"83",  x"f0",  x"af",  x"32",  x"81", -- 0D10
         x"b7",  x"cd",  x"c6",  x"f6",  x"18",  x"e0",  x"e5",  x"cd", -- 0D18
         x"97",  x"ed",  x"28",  x"ee",  x"1e",  x"24",  x"c3",  x"56", -- 0D20
         x"c3",  x"cd",  x"be",  x"c8",  x"28",  x"10",  x"cd",  x"3a", -- 0D28
         x"cd",  x"e5",  x"cd",  x"54",  x"ed",  x"cd",  x"83",  x"f0", -- 0D30
         x"cd",  x"c9",  x"e4",  x"08",  x"18",  x"c0",  x"e5",  x"11", -- 0D38
         x"5d",  x"ed",  x"18",  x"f1",  x"cd",  x"3a",  x"cd",  x"e5", -- 0D40
         x"cd",  x"54",  x"ed",  x"cd",  x"83",  x"f0",  x"cd",  x"c9", -- 0D48
         x"e4",  x"09",  x"18",  x"aa",  x"3e",  x"08",  x"f5",  x"cd", -- 0D50
         x"3f",  x"d3",  x"eb",  x"d1",  x"06",  x"00",  x"79",  x"ba", -- 0D58
         x"38",  x"01",  x"4a",  x"11",  x"ea",  x"03",  x"d5",  x"ed", -- 0D60
         x"b0",  x"af",  x"12",  x"d1",  x"c9",  x"57",  x"68",  x"e5", -- 0D68
         x"cd",  x"02",  x"f1",  x"dd",  x"cb",  x"04",  x"bf",  x"d3", -- 0D70
         x"86",  x"45",  x"21",  x"81",  x"ed",  x"e5",  x"c3",  x"20", -- 0D78
         x"c0",  x"e1",  x"16",  x"00",  x"cd",  x"02",  x"f1",  x"c3", -- 0D80
         x"8f",  x"fb",  x"cd",  x"8f",  x"fb",  x"c3",  x"cd",  x"d2", -- 0D88
         x"cd",  x"97",  x"ed",  x"07",  x"07",  x"07",  x"c9",  x"dd", -- 0D90
         x"7e",  x"08",  x"e6",  x"1c",  x"c9",  x"03",  x"92",  x"05", -- 0D98
         x"e0",  x"cf",  x"7f",  x"97",  x"c0",  x"93",  x"02",  x"cf", -- 0DA0
         x"00",  x"90",  x"01",  x"80",  x"f5",  x"e5",  x"cd",  x"6a", -- 0DA8
         x"e4",  x"e1",  x"f1",  x"ed",  x"4d",  x"ba",  x"e1",  x"57", -- 0DB0
         x"f9",  x"5c",  x"f9",  x"61",  x"f9",  x"66",  x"f9",  x"ec", -- 0DB8
         x"f0",  x"f4",  x"f0",  x"7e",  x"f9",  x"be",  x"e2",  x"87", -- 0DC0
         x"f9",  x"8f",  x"f9",  x"a5",  x"f9",  x"ac",  x"f9",  x"0d", -- 0DC8
         x"f1",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0DF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"47", -- 0DF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0E00
         x"30",  x"78",  x"78",  x"30",  x"30",  x"00",  x"30",  x"00", -- 0E08
         x"ee",  x"66",  x"cc",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0E10
         x"36",  x"36",  x"fe",  x"6c",  x"fe",  x"d8",  x"d8",  x"00", -- 0E18
         x"30",  x"7c",  x"d0",  x"7c",  x"36",  x"fc",  x"30",  x"00", -- 0E20
         x"00",  x"c6",  x"cc",  x"18",  x"30",  x"66",  x"c6",  x"00", -- 0E28
         x"38",  x"6c",  x"38",  x"76",  x"dc",  x"cc",  x"76",  x"00", -- 0E30
         x"1c",  x"0c",  x"18",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0E38
         x"18",  x"30",  x"60",  x"60",  x"60",  x"30",  x"18",  x"00", -- 0E40
         x"60",  x"30",  x"18",  x"18",  x"18",  x"30",  x"60",  x"00", -- 0E48
         x"00",  x"66",  x"3c",  x"ff",  x"3c",  x"66",  x"00",  x"00", -- 0E50
         x"00",  x"30",  x"30",  x"fc",  x"30",  x"30",  x"00",  x"00", -- 0E58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"1c",  x"0c",  x"18", -- 0E60
         x"00",  x"00",  x"00",  x"fe",  x"00",  x"00",  x"00",  x"00", -- 0E68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"30",  x"30",  x"00", -- 0E70
         x"06",  x"0c",  x"18",  x"30",  x"60",  x"c0",  x"80",  x"00", -- 0E78
         x"7c",  x"c6",  x"ce",  x"de",  x"f6",  x"e6",  x"7c",  x"00", -- 0E80
         x"30",  x"70",  x"30",  x"30",  x"30",  x"30",  x"fc",  x"00", -- 0E88
         x"78",  x"cc",  x"0c",  x"38",  x"60",  x"cc",  x"fc",  x"00", -- 0E90
         x"fc",  x"18",  x"30",  x"78",  x"0c",  x"cc",  x"78",  x"00", -- 0E98
         x"1c",  x"3c",  x"6c",  x"cc",  x"fe",  x"0c",  x"1e",  x"00", -- 0EA0
         x"fc",  x"c0",  x"f8",  x"0c",  x"0c",  x"cc",  x"78",  x"00", -- 0EA8
         x"38",  x"60",  x"c0",  x"f8",  x"cc",  x"cc",  x"78",  x"00", -- 0EB0
         x"fc",  x"cc",  x"0c",  x"18",  x"30",  x"30",  x"30",  x"00", -- 0EB8
         x"78",  x"cc",  x"cc",  x"78",  x"cc",  x"cc",  x"78",  x"00", -- 0EC0
         x"78",  x"cc",  x"cc",  x"7c",  x"0c",  x"18",  x"70",  x"00", -- 0EC8
         x"00",  x"00",  x"30",  x"30",  x"00",  x"30",  x"30",  x"00", -- 0ED0
         x"00",  x"00",  x"30",  x"30",  x"00",  x"30",  x"30",  x"60", -- 0ED8
         x"18",  x"30",  x"60",  x"c0",  x"60",  x"30",  x"18",  x"00", -- 0EE0
         x"00",  x"00",  x"fc",  x"00",  x"fc",  x"00",  x"00",  x"00", -- 0EE8
         x"60",  x"30",  x"18",  x"0c",  x"18",  x"30",  x"60",  x"00", -- 0EF0
         x"78",  x"cc",  x"0c",  x"18",  x"30",  x"00",  x"30",  x"00", -- 0EF8
         x"7c",  x"c6",  x"de",  x"d6",  x"de",  x"c0",  x"78",  x"00", -- 0F00
         x"30",  x"78",  x"cc",  x"cc",  x"fc",  x"cc",  x"cc",  x"00", -- 0F08
         x"fc",  x"66",  x"66",  x"7c",  x"66",  x"66",  x"fc",  x"00", -- 0F10
         x"3c",  x"66",  x"c0",  x"c0",  x"c0",  x"66",  x"3c",  x"00", -- 0F18
         x"f8",  x"6c",  x"66",  x"66",  x"66",  x"6c",  x"f8",  x"00", -- 0F20
         x"fe",  x"62",  x"68",  x"78",  x"68",  x"62",  x"fe",  x"00", -- 0F28
         x"fe",  x"62",  x"68",  x"78",  x"68",  x"60",  x"f0",  x"00", -- 0F30
         x"3c",  x"66",  x"c0",  x"c0",  x"ce",  x"66",  x"3c",  x"00", -- 0F38
         x"cc",  x"cc",  x"cc",  x"fc",  x"cc",  x"cc",  x"cc",  x"00", -- 0F40
         x"78",  x"30",  x"30",  x"30",  x"30",  x"30",  x"78",  x"00", -- 0F48
         x"1e",  x"0c",  x"0c",  x"0c",  x"cc",  x"cc",  x"78",  x"00", -- 0F50
         x"e6",  x"66",  x"6c",  x"70",  x"6c",  x"66",  x"e6",  x"00", -- 0F58
         x"f0",  x"60",  x"60",  x"60",  x"62",  x"66",  x"fe",  x"00", -- 0F60
         x"c6",  x"ee",  x"fe",  x"d6",  x"c6",  x"c6",  x"c6",  x"00", -- 0F68
         x"c6",  x"e6",  x"f6",  x"de",  x"ce",  x"c6",  x"c6",  x"00", -- 0F70
         x"38",  x"6c",  x"c6",  x"c6",  x"c6",  x"6c",  x"38",  x"00", -- 0F78
         x"fc",  x"66",  x"66",  x"7c",  x"60",  x"60",  x"f0",  x"00", -- 0F80
         x"78",  x"cc",  x"cc",  x"cc",  x"dc",  x"78",  x"1c",  x"00", -- 0F88
         x"fc",  x"66",  x"66",  x"7c",  x"6c",  x"66",  x"e6",  x"00", -- 0F90
         x"7c",  x"c6",  x"f0",  x"3c",  x"0e",  x"c6",  x"7c",  x"00", -- 0F98
         x"fc",  x"b4",  x"30",  x"30",  x"30",  x"30",  x"78",  x"00", -- 0FA0
         x"cc",  x"cc",  x"cc",  x"cc",  x"cc",  x"cc",  x"78",  x"00", -- 0FA8
         x"cc",  x"cc",  x"cc",  x"78",  x"78",  x"30",  x"30",  x"00", -- 0FB0
         x"c6",  x"c6",  x"c6",  x"d6",  x"fe",  x"ee",  x"c6",  x"00", -- 0FB8
         x"c6",  x"c6",  x"6c",  x"38",  x"6c",  x"c6",  x"c6",  x"00", -- 0FC0
         x"cc",  x"cc",  x"cc",  x"78",  x"30",  x"30",  x"78",  x"00", -- 0FC8
         x"fe",  x"c6",  x"8c",  x"18",  x"32",  x"66",  x"fe",  x"00", -- 0FD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0FD8
         x"18",  x"18",  x"18",  x"18",  x"18",  x"18",  x"18",  x"00", -- 0FE0
         x"00",  x"fe",  x"06",  x"06",  x"00",  x"00",  x"00",  x"00", -- 0FE8
         x"10",  x"38",  x"6c",  x"c6",  x"00",  x"00",  x"00",  x"00", -- 0FF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"ff", -- 0FF8
         x"c3",  x"5f",  x"f1",  x"18",  x"4c",  x"00",  x"18",  x"67", -- 1000
         x"02",  x"18",  x"62",  x"03",  x"18",  x"2b",  x"04",  x"c3", -- 1008
         x"b7",  x"f0",  x"c3",  x"66",  x"f1",  x"c3",  x"2d",  x"f0", -- 1010
         x"c3",  x"83",  x"f0",  x"c3",  x"a0",  x"f0",  x"c3",  x"24", -- 1018
         x"f0",  x"c3",  x"c9",  x"e4",  x"c5",  x"cd",  x"83",  x"f0", -- 1020
         x"cd",  x"6f",  x"f0",  x"18",  x"07",  x"c5",  x"cd",  x"83", -- 1028
         x"f0",  x"cd",  x"6d",  x"f0",  x"cd",  x"a0",  x"f0",  x"c1", -- 1030
         x"c9",  x"cd",  x"48",  x"f0",  x"cd",  x"6d",  x"f0",  x"f5", -- 1038
         x"db",  x"88",  x"e6",  x"fb",  x"d3",  x"88",  x"f1",  x"c9", -- 1040
         x"f5",  x"db",  x"88",  x"f6",  x"04",  x"d3",  x"88",  x"f1", -- 1048
         x"c9",  x"f3",  x"e5",  x"e1",  x"e1",  x"23",  x"e5",  x"2b", -- 1050
         x"3b",  x"3b",  x"fb",  x"f5",  x"d5",  x"5e",  x"16",  x"00", -- 1058
         x"2a",  x"b0",  x"b7",  x"19",  x"19",  x"5e",  x"23",  x"56", -- 1060
         x"eb",  x"d1",  x"f1",  x"e3",  x"c9",  x"37",  x"ed",  x"a7", -- 1068
         x"e5",  x"d5",  x"c5",  x"e5",  x"21",  x"ec",  x"f3",  x"e3", -- 1070
         x"e5",  x"f5",  x"d5",  x"38",  x"e1",  x"3a",  x"80",  x"b7", -- 1078
         x"5f",  x"18",  x"db",  x"c1",  x"fd",  x"e5",  x"fd",  x"21", -- 1080
         x"00",  x"00",  x"fd",  x"39",  x"f3",  x"dd",  x"77",  x"0b", -- 1088
         x"db",  x"88",  x"f6",  x"24",  x"d3",  x"88",  x"ed",  x"7b", -- 1090
         x"ae",  x"b7",  x"fb",  x"dd",  x"7e",  x"0b",  x"c5",  x"c9", -- 1098
         x"c1",  x"dd",  x"77",  x"0b",  x"db",  x"88",  x"cb",  x"97", -- 10A0
         x"cb",  x"af",  x"f3",  x"d3",  x"88",  x"fd",  x"f9",  x"fb", -- 10A8
         x"dd",  x"7e",  x"0b",  x"fd",  x"e1",  x"c5",  x"c9",  x"e3", -- 10B0
         x"d5",  x"5e",  x"23",  x"56",  x"23",  x"eb",  x"19",  x"e3", -- 10B8
         x"eb",  x"f3",  x"33",  x"33",  x"e3",  x"3b",  x"3b",  x"fb", -- 10C0
         x"c9",  x"dd",  x"7e",  x"02",  x"cd",  x"c4",  x"f3",  x"e3", -- 10C8
         x"cd",  x"06",  x"f9",  x"e3",  x"c9",  x"7f",  x"7f",  x"53", -- 10D0
         x"57",  x"49",  x"54",  x"43",  x"48",  x"01",  x"a7",  x"28", -- 10D8
         x"08",  x"cd",  x"8f",  x"fb",  x"cd",  x"31",  x"c3",  x"18", -- 10E0
         x"21",  x"cd",  x"f4",  x"f0",  x"cd",  x"8f",  x"fb",  x"cd", -- 10E8
         x"75",  x"c2",  x"18",  x"06",  x"cd",  x"8f",  x"fb",  x"cd", -- 10F0
         x"a1",  x"c1",  x"ed",  x"5b",  x"a0",  x"b7",  x"18",  x"0a", -- 10F8
         x"2e",  x"02",  x"3e",  x"02",  x"cd",  x"8f",  x"fb",  x"cd", -- 1100
         x"9c",  x"c3",  x"c3",  x"9c",  x"fb",  x"cd",  x"8f",  x"fb", -- 1108
         x"cd",  x"56",  x"d6",  x"18",  x"e5",  x"7f",  x"7f",  x"4a", -- 1110
         x"55",  x"4d",  x"50",  x"03",  x"7d",  x"b7",  x"28",  x"46", -- 1118
         x"47",  x"0e",  x"80",  x"ed",  x"78",  x"3c",  x"20",  x"13", -- 1120
         x"cd",  x"cf",  x"f0",  x"4b",  x"65",  x"69",  x"6e",  x"20", -- 1128
         x"4d",  x"6f",  x"64",  x"75",  x"6c",  x"21",  x"07",  x"0d", -- 1130
         x"0a",  x"00",  x"c9",  x"c5",  x"26",  x"b8",  x"06",  x"07", -- 1138
         x"04",  x"28",  x"0d",  x"ed",  x"78",  x"2f",  x"e6",  x"70", -- 1140
         x"20",  x"f6",  x"ed",  x"79",  x"68",  x"77",  x"18",  x"f0", -- 1148
         x"c1",  x"3e",  x"fd",  x"68",  x"77",  x"f3",  x"ed",  x"79", -- 1150
         x"db",  x"88",  x"e6",  x"7e",  x"c3",  x"b4",  x"b7",  x"3e", -- 1158
         x"e3",  x"d3",  x"86",  x"c3",  x"51",  x"c0",  x"31",  x"c4", -- 1160
         x"01",  x"3e",  x"e3",  x"d3",  x"86",  x"cd",  x"91",  x"c0", -- 1168
         x"cd",  x"f0",  x"c9",  x"cd",  x"9c",  x"fb",  x"01",  x"80", -- 1170
         x"08",  x"ed",  x"78",  x"3d",  x"20",  x"14",  x"3e",  x"41", -- 1178
         x"ed",  x"79",  x"32",  x"08",  x"b8",  x"dd",  x"7e",  x"04", -- 1180
         x"e6",  x"fc",  x"dd",  x"77",  x"04",  x"d3",  x"86",  x"c3", -- 1188
         x"00",  x"40",  x"06",  x"fc",  x"ed",  x"78",  x"fe",  x"a7", -- 1190
         x"20",  x"37",  x"01",  x"f3",  x"b3",  x"ed",  x"78",  x"3d", -- 1198
         x"28",  x"2f",  x"fe",  x"04",  x"28",  x"2b",  x"cd",  x"cf", -- 11A0
         x"f0",  x"0c",  x"0a",  x"41",  x"75",  x"74",  x"6f",  x"73", -- 11A8
         x"74",  x"61",  x"72",  x"74",  x"20",  x"46",  x"6c",  x"6f", -- 11B0
         x"70",  x"70",  x"79",  x"0d",  x"0a",  x"00",  x"06",  x"00", -- 11B8
         x"cd",  x"7c",  x"e3",  x"38",  x"0c",  x"10",  x"f9",  x"3e", -- 11C0
         x"01",  x"32",  x"81",  x"b7",  x"3e",  x"fc",  x"cd",  x"1d", -- 11C8
         x"f1",  x"af",  x"32",  x"81",  x"b7",  x"18",  x"08",  x"7f", -- 11D0
         x"7f",  x"4d",  x"45",  x"4e",  x"55",  x"01",  x"e1",  x"cd", -- 11D8
         x"cf",  x"f0",  x"0c",  x"0a",  x"2a",  x"20",  x"4b",  x"43", -- 11E0
         x"2d",  x"43",  x"41",  x"4f",  x"53",  x"20",  x"34",  x"2e", -- 11E8
         x"37",  x"20",  x"00",  x"cd",  x"d2",  x"fb",  x"cd",  x"cf", -- 11F0
         x"f0",  x"20",  x"2a",  x"00",  x"2a",  x"81",  x"b7",  x"1e", -- 11F8
         x"00",  x"2d",  x"20",  x"01",  x"5c",  x"21",  x"00",  x"c0", -- 1200
         x"4d",  x"45",  x"cd",  x"db",  x"f4",  x"3e",  x"02",  x"cd", -- 1208
         x"a6",  x"f3",  x"cd",  x"7c",  x"e3",  x"38",  x"62",  x"dd", -- 1210
         x"7e",  x"09",  x"ed",  x"b1",  x"e2",  x"79",  x"f2",  x"ed", -- 1218
         x"a1",  x"e2",  x"79",  x"f2",  x"20",  x"f4",  x"7e",  x"fe", -- 1220
         x"20",  x"38",  x"27",  x"cb",  x"43",  x"28",  x"06",  x"fe", -- 1228
         x"7b",  x"30",  x"da",  x"18",  x"10",  x"fe",  x"30",  x"38", -- 1230
         x"d4",  x"fe",  x"5b",  x"30",  x"d0",  x"fe",  x"41",  x"30", -- 1238
         x"04",  x"fe",  x"3b",  x"30",  x"c8",  x"cd",  x"d5",  x"f3", -- 1240
         x"23",  x"0b",  x"79",  x"b0",  x"20",  x"d8",  x"3e",  x"02", -- 1248
         x"18",  x"24",  x"cb",  x"4b",  x"28",  x"b4",  x"3a",  x"9e", -- 1250
         x"b7",  x"fe",  x"0f",  x"38",  x"ad",  x"3e",  x"0b",  x"32", -- 1258
         x"a0",  x"b7",  x"23",  x"cd",  x"b4",  x"f3",  x"2b",  x"18", -- 1260
         x"a1",  x"db",  x"88",  x"e6",  x"df",  x"f6",  x"04",  x"d3", -- 1268
         x"88",  x"cd",  x"9c",  x"fb",  x"3e",  x"0d",  x"cd",  x"a6", -- 1270
         x"f3",  x"cd",  x"7e",  x"f2",  x"18",  x"eb",  x"cd",  x"99", -- 1278
         x"f4",  x"30",  x"0a",  x"3e",  x"0b",  x"cd",  x"8c",  x"e0", -- 1280
         x"3e",  x"02",  x"c3",  x"8c",  x"e0",  x"13",  x"1a",  x"e6", -- 1288
         x"df",  x"c8",  x"3a",  x"02",  x"b8",  x"32",  x"80",  x"b7", -- 1290
         x"cd",  x"51",  x"f3",  x"38",  x"3f",  x"3a",  x"05",  x"b8", -- 1298
         x"e6",  x"01",  x"20",  x"0a",  x"cd",  x"8f",  x"fb",  x"06", -- 12A0
         x"20",  x"cd",  x"53",  x"f3",  x"38",  x"2e",  x"d5",  x"16", -- 12A8
         x"d1",  x"cd",  x"00",  x"f1",  x"dd",  x"cb",  x"04",  x"bf", -- 12B0
         x"d3",  x"86",  x"eb",  x"e3",  x"eb",  x"06",  x"20",  x"cd", -- 12B8
         x"53",  x"f3",  x"38",  x"13",  x"eb",  x"e3",  x"eb",  x"3e", -- 12C0
         x"10",  x"82",  x"57",  x"30",  x"e4",  x"ed",  x"5b",  x"7f", -- 12C8
         x"b7",  x"cd",  x"00",  x"f1",  x"d1",  x"18",  x"2c",  x"f1", -- 12D0
         x"af",  x"32",  x"05",  x"b8",  x"7e",  x"23",  x"e5",  x"fe", -- 12D8
         x"1f",  x"c8",  x"f5",  x"cd",  x"20",  x"f5",  x"c1",  x"38", -- 12E0
         x"46",  x"3a",  x"81",  x"b7",  x"48",  x"cb",  x"a0",  x"cb", -- 12E8
         x"28",  x"b8",  x"38",  x"2d",  x"28",  x"04",  x"cb",  x"61", -- 12F0
         x"20",  x"19",  x"cb",  x"41",  x"cd",  x"ff",  x"f5",  x"c0", -- 12F8
         x"c3",  x"3f",  x"f0",  x"cd",  x"cf",  x"f0",  x"4b",  x"6f", -- 1300
         x"6d",  x"6d",  x"61",  x"6e",  x"64",  x"6f",  x"3f",  x"07", -- 1308
         x"00",  x"18",  x"3b",  x"cd",  x"cf",  x"f0",  x"5a",  x"75", -- 1310
         x"20",  x"76",  x"69",  x"65",  x"6c",  x"65",  x"00",  x"18", -- 1318
         x"1d",  x"cd",  x"cf",  x"f0",  x"5a",  x"75",  x"20",  x"77", -- 1320
         x"65",  x"6e",  x"69",  x"67",  x"00",  x"18",  x"0f",  x"cd", -- 1328
         x"cf",  x"f0",  x"46",  x"65",  x"68",  x"6c",  x"65",  x"72", -- 1330
         x"68",  x"61",  x"66",  x"74",  x"65",  x"00",  x"e1",  x"cd", -- 1338
         x"cf",  x"f0",  x"20",  x"41",  x"72",  x"67",  x"75",  x"6d", -- 1340
         x"65",  x"6e",  x"74",  x"65",  x"07",  x"00",  x"c3",  x"db", -- 1348
         x"f4",  x"06",  x"00",  x"21",  x"00",  x"c0",  x"4d",  x"dd", -- 1350
         x"7e",  x"09",  x"ed",  x"b1",  x"37",  x"3f",  x"e0",  x"ed", -- 1358
         x"a1",  x"20",  x"f7",  x"f5",  x"d5",  x"1a",  x"13",  x"fe", -- 1360
         x"21",  x"38",  x"0d",  x"cb",  x"6e",  x"cc",  x"3d",  x"f5", -- 1368
         x"ed",  x"a1",  x"28",  x"f1",  x"d1",  x"f1",  x"18",  x"e2", -- 1370
         x"7e",  x"fe",  x"20",  x"38",  x"08",  x"fe",  x"80",  x"30", -- 1378
         x"f3",  x"23",  x"0b",  x"18",  x"f3",  x"f1",  x"f1",  x"37", -- 1380
         x"c9",  x"cd",  x"99",  x"f3",  x"21",  x"05",  x"f0",  x"e5", -- 1388
         x"2a",  x"b9",  x"b7",  x"e3",  x"22",  x"b9",  x"b7",  x"e1", -- 1390
         x"c9",  x"21",  x"0e",  x"f0",  x"e5",  x"2a",  x"bb",  x"b7", -- 1398
         x"e3",  x"22",  x"bb",  x"b7",  x"e1",  x"c9",  x"cd",  x"8c", -- 13A0
         x"e0",  x"3a",  x"ec",  x"b7",  x"fe",  x"20",  x"30",  x"02", -- 13A8
         x"3e",  x"25",  x"18",  x"21",  x"7c",  x"cd",  x"c4",  x"f3", -- 13B0
         x"7d",  x"cd",  x"c4",  x"f3",  x"3e",  x"20",  x"18",  x"15", -- 13B8
         x"3e",  x"10",  x"18",  x"11",  x"f5",  x"0f",  x"0f",  x"0f", -- 13C0
         x"0f",  x"cd",  x"cd",  x"f3",  x"f1",  x"e6",  x"0f",  x"c6", -- 13C8
         x"90",  x"27",  x"ce",  x"40",  x"27",  x"e5",  x"2a",  x"b9", -- 13D0
         x"b7",  x"d5",  x"c5",  x"5e",  x"16",  x"00",  x"2a",  x"b0", -- 13D8
         x"b7",  x"f5",  x"19",  x"19",  x"f1",  x"5e",  x"23",  x"56", -- 13E0
         x"eb",  x"cd",  x"b9",  x"e1",  x"c1",  x"d1",  x"e1",  x"c9", -- 13E8
         x"e5",  x"2a",  x"bb",  x"b7",  x"18",  x"e3",  x"e5",  x"d5", -- 13F0
         x"c5",  x"dd",  x"cb",  x"08",  x"76",  x"20",  x"60",  x"1e", -- 13F8
         x"00",  x"cd",  x"51",  x"f0",  x"25",  x"1c",  x"06",  x"0f", -- 1400
         x"cd",  x"73",  x"e3",  x"38",  x"07",  x"0b",  x"78",  x"b1", -- 1408
         x"20",  x"f6",  x"18",  x"ed",  x"cb",  x"43",  x"28",  x"04", -- 1410
         x"cd",  x"51",  x"f0",  x"25",  x"57",  x"dd",  x"cb",  x"08", -- 1418
         x"6e",  x"c4",  x"b1",  x"e2",  x"7a",  x"21",  x"a2",  x"b7", -- 1420
         x"cb",  x"66",  x"28",  x"0d",  x"ed",  x"5b",  x"a0",  x"b7", -- 1428
         x"cd",  x"83",  x"e1",  x"ed",  x"53",  x"a0",  x"b7",  x"18", -- 1430
         x"c6",  x"fe",  x"1b",  x"20",  x"04",  x"cb",  x"e6",  x"18", -- 1438
         x"be",  x"fe",  x"f1",  x"38",  x"a7",  x"e6",  x"0f",  x"47", -- 1440
         x"21",  x"00",  x"b9",  x"7e",  x"2c",  x"28",  x"b0",  x"a7", -- 1448
         x"20",  x"f9",  x"10",  x"f7",  x"7d",  x"fe",  x"9c",  x"30", -- 1450
         x"a6",  x"dd",  x"cb",  x"08",  x"f6",  x"18",  x"08",  x"cd", -- 1458
         x"7c",  x"e3",  x"38",  x"1a",  x"2a",  x"d1",  x"b7",  x"7e", -- 1460
         x"fe",  x"1b",  x"20",  x"0b",  x"23",  x"22",  x"d1",  x"b7", -- 1468
         x"21",  x"a2",  x"b7",  x"cb",  x"e6",  x"18",  x"82",  x"23", -- 1470
         x"22",  x"d1",  x"b7",  x"a7",  x"20",  x"06",  x"dd",  x"cb", -- 1478
         x"08",  x"b6",  x"18",  x"bb",  x"21",  x"a2",  x"b7",  x"cb", -- 1480
         x"66",  x"ca",  x"ec",  x"f3",  x"ed",  x"5b",  x"a0",  x"b7", -- 1488
         x"cd",  x"83",  x"e1",  x"ed",  x"53",  x"a0",  x"b7",  x"18", -- 1490
         x"dc",  x"cd",  x"f0",  x"f3",  x"cd",  x"d5",  x"f3",  x"fe", -- 1498
         x"03",  x"37",  x"28",  x"04",  x"fe",  x"0d",  x"20",  x"f1", -- 14A0
         x"f5",  x"cd",  x"db",  x"f4",  x"ed",  x"5b",  x"a0",  x"b7", -- 14A8
         x"ba",  x"20",  x"04",  x"3a",  x"9f",  x"b7",  x"57",  x"15", -- 14B0
         x"e5",  x"cd",  x"68",  x"e0",  x"eb",  x"e1",  x"f1",  x"c9", -- 14B8
         x"7f",  x"7f",  x"67",  x"6f",  x"03",  x"e5",  x"eb",  x"50", -- 14C0
         x"59",  x"ed",  x"4b",  x"88",  x"b7",  x"3a",  x"8a",  x"b7", -- 14C8
         x"c9",  x"cd",  x"cf",  x"f0",  x"45",  x"52",  x"52",  x"4f", -- 14D0
         x"52",  x"07",  x"00",  x"cd",  x"cf",  x"f0",  x"0d",  x"0a", -- 14D8
         x"00",  x"c9",  x"cd",  x"e5",  x"f4",  x"cd",  x"b4",  x"f3", -- 14E0
         x"eb",  x"c9",  x"13",  x"1a",  x"fe",  x"20",  x"28",  x"fa", -- 14E8
         x"af",  x"21",  x"98",  x"b7",  x"77",  x"2b",  x"77",  x"2b", -- 14F0
         x"77",  x"1a",  x"b7",  x"c8",  x"fe",  x"20",  x"c8",  x"d6", -- 14F8
         x"30",  x"d8",  x"fe",  x"0a",  x"38",  x"0b",  x"d6",  x"07", -- 1500
         x"e6",  x"df",  x"fe",  x"0a",  x"d8",  x"fe",  x"10",  x"3f", -- 1508
         x"d8",  x"13",  x"34",  x"23",  x"ed",  x"6f",  x"23",  x"ed", -- 1510
         x"6f",  x"2b",  x"2b",  x"28",  x"dc",  x"1b",  x"37",  x"c9", -- 1518
         x"01",  x"81",  x"b7",  x"af",  x"02",  x"cd",  x"eb",  x"f4", -- 1520
         x"d8",  x"7e",  x"b7",  x"c8",  x"23",  x"03",  x"7e",  x"02", -- 1528
         x"23",  x"03",  x"7e",  x"02",  x"2e",  x"81",  x"34",  x"7e", -- 1530
         x"c6",  x"f5",  x"30",  x"e9",  x"c9",  x"fe",  x"61",  x"d8", -- 1538
         x"fe",  x"7b",  x"d0",  x"e6",  x"df",  x"c9",  x"dd",  x"36", -- 1540
         x"05",  x"00",  x"dd",  x"36",  x"06",  x"b7",  x"c9",  x"c5", -- 1548
         x"4e",  x"23",  x"46",  x"23",  x"ed",  x"b3",  x"c1",  x"c9", -- 1550
         x"56",  x"23",  x"cd",  x"4f",  x"f5",  x"15",  x"20",  x"fa", -- 1558
         x"c9",  x"f3",  x"cd",  x"5a",  x"f5",  x"fb",  x"c9",  x"21", -- 1560
         x"06",  x"00",  x"cd",  x"cf",  x"f0",  x"4e",  x"61",  x"6d", -- 1568
         x"65",  x"20",  x"3a",  x"00",  x"cd",  x"99",  x"f4",  x"d8", -- 1570
         x"19",  x"c9",  x"7f",  x"7f",  x"53",  x"41",  x"56",  x"45", -- 1578
         x"05",  x"cd",  x"67",  x"f5",  x"d8",  x"cd",  x"c0",  x"e4", -- 1580
         x"e5",  x"01",  x"0b",  x"00",  x"ed",  x"b0",  x"af",  x"12", -- 1588
         x"21",  x"81",  x"b7",  x"1e",  x"10",  x"0e",  x"15",  x"ed", -- 1590
         x"b0",  x"cd",  x"46",  x"f5",  x"e1",  x"cd",  x"c9",  x"e4", -- 1598
         x"02",  x"d8",  x"2a",  x"84",  x"b7",  x"ed",  x"5b",  x"82", -- 15A0
         x"b7",  x"a7",  x"ed",  x"52",  x"e5",  x"2a",  x"82",  x"b7", -- 15A8
         x"11",  x"00",  x"b7",  x"01",  x"80",  x"00",  x"3a",  x"01", -- 15B0
         x"b8",  x"e6",  x"01",  x"20",  x"0f",  x"41",  x"cd",  x"3f", -- 15B8
         x"f0",  x"7e",  x"cd",  x"48",  x"f0",  x"12",  x"23",  x"13", -- 15C0
         x"10",  x"f4",  x"18",  x"02",  x"ed",  x"b0",  x"22",  x"82", -- 15C8
         x"b7",  x"e1",  x"cd",  x"cf",  x"f0",  x"02",  x"00",  x"cd", -- 15D0
         x"c9",  x"f0",  x"00",  x"cd",  x"7c",  x"e3",  x"01",  x"a0", -- 15D8
         x"00",  x"38",  x"11",  x"11",  x"80",  x"00",  x"ed",  x"52", -- 15E0
         x"28",  x"0a",  x"38",  x"08",  x"e5",  x"cd",  x"c9",  x"e4", -- 15E8
         x"00",  x"30",  x"ba",  x"e1",  x"cd",  x"c9",  x"e4",  x"03", -- 15F0
         x"cd",  x"c0",  x"e4",  x"cd",  x"db",  x"f4",  x"c9",  x"ed", -- 15F8
         x"4b",  x"86",  x"b7",  x"ed",  x"5b",  x"84",  x"b7",  x"2a", -- 1600
         x"82",  x"b7",  x"3a",  x"81",  x"b7",  x"c9",  x"dd",  x"34", -- 1608
         x"03",  x"cd",  x"c9",  x"e4",  x"01",  x"30",  x"25",  x"cd", -- 1610
         x"97",  x"ed",  x"37",  x"c0",  x"cd",  x"cf",  x"f0",  x"09", -- 1618
         x"09",  x"09",  x"20",  x"00",  x"cd",  x"c9",  x"f0",  x"20", -- 1620
         x"3f",  x"1e",  x"00",  x"dd",  x"7e",  x"03",  x"3d",  x"28", -- 1628
         x"e0",  x"cd",  x"f6",  x"f3",  x"fe",  x"03",  x"37",  x"c8", -- 1630
         x"fe",  x"0a",  x"20",  x"d5",  x"dd",  x"7e",  x"02",  x"dd", -- 1638
         x"46",  x"03",  x"05",  x"28",  x"17",  x"04",  x"b8",  x"28", -- 1640
         x"0b",  x"3c",  x"28",  x"08",  x"cd",  x"c9",  x"f0",  x"2a", -- 1648
         x"19",  x"00",  x"18",  x"bd",  x"cd",  x"c9",  x"f0",  x"3e", -- 1650
         x"20",  x"19",  x"00",  x"c9",  x"3d",  x"20",  x"ed",  x"21", -- 1658
         x"00",  x"b7",  x"06",  x"0b",  x"7e",  x"b7",  x"28",  x"10", -- 1660
         x"fe",  x"20",  x"38",  x"20",  x"fe",  x"7f",  x"38",  x"08", -- 1668
         x"fe",  x"d3",  x"38",  x"18",  x"fe",  x"d6",  x"30",  x"14", -- 1670
         x"2c",  x"10",  x"e9",  x"2e",  x"00",  x"06",  x"0b",  x"7e", -- 1678
         x"e6",  x"7f",  x"23",  x"b7",  x"c4",  x"8c",  x"e0",  x"10", -- 1680
         x"f6",  x"cd",  x"bc",  x"f3",  x"a7",  x"c9",  x"cd",  x"cf", -- 1688
         x"f0",  x"4b",  x"65",  x"69",  x"6e",  x"65",  x"20",  x"4d", -- 1690
         x"43",  x"2d",  x"44",  x"61",  x"74",  x"65",  x"69",  x"21", -- 1698
         x"00",  x"cd",  x"8f",  x"e5",  x"37",  x"c9",  x"7f",  x"7f", -- 16A0
         x"56",  x"45",  x"52",  x"49",  x"46",  x"59",  x"01",  x"cd", -- 16A8
         x"97",  x"ed",  x"c0",  x"dd",  x"77",  x"07",  x"18",  x"1d", -- 16B0
         x"7f",  x"7f",  x"4c",  x"4f",  x"41",  x"44",  x"01",  x"cd", -- 16B8
         x"97",  x"ed",  x"c4",  x"67",  x"f5",  x"d8",  x"dd",  x"36", -- 16C0
         x"07",  x"01",  x"3a",  x"81",  x"b7",  x"fe",  x"02",  x"38", -- 16C8
         x"04",  x"dd",  x"cb",  x"07",  x"ce",  x"cd",  x"46",  x"f5", -- 16D0
         x"cd",  x"c9",  x"e4",  x"04",  x"30",  x"05",  x"cd",  x"97", -- 16D8
         x"ed",  x"37",  x"c0",  x"cd",  x"15",  x"f6",  x"38",  x"b9", -- 16E0
         x"dd",  x"cb",  x"07",  x"46",  x"28",  x"4d",  x"2e",  x"10", -- 16E8
         x"7e",  x"07",  x"07",  x"dd",  x"ae",  x"07",  x"e6",  x"1c", -- 16F0
         x"dd",  x"ae",  x"07",  x"dd",  x"77",  x"07",  x"7e",  x"d6", -- 16F8
         x"02",  x"fe",  x"09",  x"30",  x"89",  x"2a",  x"15",  x"b7", -- 1700
         x"e5",  x"ed",  x"5b",  x"13",  x"b7",  x"2a",  x"11",  x"b7", -- 1708
         x"3a",  x"81",  x"b7",  x"a7",  x"28",  x"11",  x"ed",  x"4b", -- 1710
         x"82",  x"b7",  x"09",  x"eb",  x"09",  x"eb",  x"dd",  x"cb", -- 1718
         x"07",  x"66",  x"20",  x"03",  x"e3",  x"09",  x"e3",  x"cd", -- 1720
         x"e2",  x"f4",  x"3a",  x"10",  x"b7",  x"fe",  x"03",  x"38", -- 1728
         x"05",  x"e3",  x"cd",  x"b4",  x"f3",  x"e3",  x"c1",  x"ed", -- 1730
         x"43",  x"86",  x"b7",  x"cd",  x"db",  x"f4",  x"eb",  x"cd", -- 1738
         x"0e",  x"f6",  x"38",  x"a2",  x"dd",  x"cb",  x"07",  x"46", -- 1740
         x"28",  x"25",  x"e5",  x"ed",  x"52",  x"01",  x"80",  x"00", -- 1748
         x"ed",  x"42",  x"09",  x"30",  x"01",  x"4d",  x"21",  x"00", -- 1750
         x"b7",  x"3a",  x"01",  x"b8",  x"e6",  x"01",  x"20",  x"16", -- 1758
         x"41",  x"7e",  x"cd",  x"3f",  x"f0",  x"12",  x"23",  x"13", -- 1760
         x"cd",  x"48",  x"f0",  x"10",  x"f4",  x"18",  x"09",  x"dd", -- 1768
         x"34",  x"02",  x"28",  x"0a",  x"18",  x"c9",  x"ed",  x"b0", -- 1770
         x"e1",  x"ed",  x"52",  x"19",  x"20",  x"c1",  x"cd",  x"c0", -- 1778
         x"e4",  x"cd",  x"db",  x"f4",  x"cd",  x"c9",  x"e4",  x"05", -- 1780
         x"d8",  x"dd",  x"7e",  x"07",  x"e6",  x"03",  x"3d",  x"c0", -- 1788
         x"dd",  x"7e",  x"07",  x"e6",  x"1c",  x"fe",  x"0c",  x"dd", -- 1790
         x"36",  x"07",  x"00",  x"3f",  x"d0",  x"2a",  x"86",  x"b7", -- 1798
         x"e9",  x"7f",  x"7f",  x"43",  x"4f",  x"4c",  x"4f",  x"52", -- 17A0
         x"01",  x"cd",  x"8f",  x"fb",  x"c3",  x"66",  x"c5",  x"cd", -- 17A8
         x"8f",  x"fb",  x"c3",  x"80",  x"c5",  x"e5",  x"21",  x"a2", -- 17B0
         x"b7",  x"cb",  x"de",  x"cd",  x"d5",  x"f3",  x"cb",  x"9e", -- 17B8
         x"e1",  x"c9",  x"7f",  x"7f",  x"44",  x"49",  x"53",  x"50", -- 17C0
         x"4c",  x"41",  x"59",  x"03",  x"cd",  x"8f",  x"fb",  x"cd", -- 17C8
         x"fd",  x"c7",  x"18",  x"0f",  x"7f",  x"7f",  x"4d",  x"4f", -- 17D0
         x"44",  x"49",  x"46",  x"59",  x"03",  x"cd",  x"8f",  x"fb", -- 17D8
         x"cd",  x"2e",  x"c8",  x"c3",  x"9c",  x"fb",  x"7f",  x"7f", -- 17E0
         x"57",  x"49",  x"4e",  x"44",  x"4f",  x"57",  x"01",  x"cd", -- 17E8
         x"8f",  x"fb",  x"cd",  x"9b",  x"c5",  x"18",  x"ec",  x"cd", -- 17F0
         x"8f",  x"fb",  x"cd",  x"fa",  x"c5",  x"18",  x"e4",  x"cd", -- 17F8
         x"8f",  x"fb",  x"cd",  x"ca",  x"c5",  x"18",  x"dc",  x"7f", -- 1800
         x"7f",  x"4b",  x"45",  x"59",  x"01",  x"fe",  x"01",  x"30", -- 1808
         x"08",  x"cd",  x"8f",  x"fb",  x"cd",  x"1c",  x"c5",  x"18", -- 1810
         x"ca",  x"7d",  x"cd",  x"8f",  x"fb",  x"cd",  x"70",  x"c4", -- 1818
         x"18",  x"c1",  x"d5",  x"f5",  x"e5",  x"cd",  x"3e",  x"e0", -- 1820
         x"38",  x"22",  x"e5",  x"cd",  x"68",  x"e0",  x"7e",  x"e1", -- 1828
         x"a7",  x"20",  x"0a",  x"3e",  x"06",  x"b5",  x"6f",  x"7e", -- 1830
         x"ee",  x"7f",  x"77",  x"18",  x"0f",  x"c5",  x"ed",  x"5b", -- 1838
         x"ee",  x"b7",  x"06",  x"08",  x"1a",  x"ae",  x"77",  x"13", -- 1840
         x"2c",  x"10",  x"f9",  x"c1",  x"e1",  x"f1",  x"d1",  x"c9", -- 1848
         x"cd",  x"8f",  x"fb",  x"cd",  x"74",  x"c7",  x"18",  x"16", -- 1850
         x"cd",  x"8f",  x"fb",  x"cd",  x"7f",  x"c7",  x"18",  x"0e", -- 1858
         x"cd",  x"8f",  x"fb",  x"cd",  x"ad",  x"c6",  x"18",  x"06", -- 1860
         x"cd",  x"8f",  x"fb",  x"cd",  x"30",  x"c6",  x"c3",  x"9c", -- 1868
         x"fb",  x"cd",  x"8f",  x"fb",  x"cd",  x"79",  x"cd",  x"18", -- 1870
         x"06",  x"cd",  x"8f",  x"fb",  x"cd",  x"e3",  x"cc",  x"cd", -- 1878
         x"9c",  x"fb",  x"d0",  x"2a",  x"c9",  x"b7",  x"cd",  x"a0", -- 1880
         x"f0",  x"e9",  x"e5",  x"c5",  x"cd",  x"83",  x"f0",  x"cb", -- 1888
         x"6b",  x"20",  x"59",  x"d5",  x"23",  x"23",  x"cb",  x"7b", -- 1890
         x"20",  x"47",  x"e5",  x"7b",  x"e6",  x"07",  x"21",  x"f0", -- 1898
         x"fd",  x"85",  x"6f",  x"7a",  x"53",  x"5e",  x"e1",  x"cd", -- 18A0
         x"6d",  x"f0",  x"d1",  x"57",  x"7b",  x"e6",  x"4f",  x"ee", -- 18A8
         x"43",  x"20",  x"25",  x"cd",  x"97",  x"ed",  x"20",  x"20", -- 18B0
         x"cd",  x"cf",  x"f0",  x"56",  x"45",  x"52",  x"49",  x"46", -- 18B8
         x"59",  x"20",  x"3f",  x"28",  x"59",  x"29",  x"3a",  x"00", -- 18C0
         x"cd",  x"f6",  x"f3",  x"cd",  x"b5",  x"f7",  x"f5",  x"cd", -- 18C8
         x"db",  x"f4",  x"f1",  x"fe",  x"59",  x"cc",  x"af",  x"f6", -- 18D0
         x"7a",  x"cb",  x"9b",  x"cd",  x"a0",  x"f0",  x"c1",  x"e1", -- 18D8
         x"c9",  x"cd",  x"68",  x"e3",  x"d1",  x"57",  x"30",  x"f0", -- 18E0
         x"cb",  x"bb",  x"18",  x"ec",  x"3a",  x"5e",  x"03",  x"a7", -- 18E8
         x"28",  x"09",  x"cd",  x"a0",  x"f0",  x"cd",  x"41",  x"c6", -- 18F0
         x"cd",  x"83",  x"f0",  x"16",  x"00",  x"cd",  x"00",  x"f1", -- 18F8
         x"c3",  x"69",  x"f2",  x"cd",  x"d5",  x"f3",  x"7e",  x"23", -- 1900
         x"a7",  x"20",  x"f8",  x"c9",  x"cd",  x"ff",  x"f5",  x"dd", -- 1908
         x"cb",  x"08",  x"4e",  x"20",  x"fa",  x"79",  x"e6",  x"1e", -- 1910
         x"ee",  x"9f",  x"4f",  x"78",  x"a7",  x"f3",  x"28",  x"0d", -- 1918
         x"cb",  x"b9",  x"dd",  x"cb",  x"08",  x"ce",  x"3e",  x"c7", -- 1920
         x"d3",  x"8e",  x"78",  x"d3",  x"8e",  x"db",  x"89",  x"e6", -- 1928
         x"60",  x"b1",  x"d3",  x"89",  x"fb",  x"0e",  x"8c",  x"cd", -- 1930
         x"3c",  x"f9",  x"0c",  x"eb",  x"7d",  x"a7",  x"2e",  x"03", -- 1938
         x"28",  x"0c",  x"6f",  x"3e",  x"38",  x"cb",  x"3c",  x"1f", -- 1940
         x"1f",  x"1f",  x"f3",  x"ed",  x"79",  x"fb",  x"ed",  x"69", -- 1948
         x"c9",  x"21",  x"a2",  x"b7",  x"cb",  x"e6",  x"c9",  x"01", -- 1950
         x"00",  x"b2",  x"18",  x"0d",  x"01",  x"05",  x"ad",  x"18", -- 1958
         x"08",  x"01",  x"04",  x"ad",  x"18",  x"03",  x"01",  x"01", -- 1960
         x"b2",  x"60",  x"2e",  x"00",  x"22",  x"cb",  x"b7",  x"06", -- 1968
         x"fa",  x"78",  x"f3",  x"dd",  x"a6",  x"01",  x"a9",  x"dd", -- 1970
         x"77",  x"01",  x"d3",  x"84",  x"fb",  x"c9",  x"0e",  x"04", -- 1978
         x"21",  x"a2",  x"b7",  x"7e",  x"a9",  x"77",  x"c9",  x"f3", -- 1980
         x"dd",  x"7e",  x"01",  x"ee",  x"02",  x"18",  x"e8",  x"21", -- 1988
         x"a2",  x"b7",  x"cb",  x"b6",  x"01",  x"08",  x"ff",  x"cd", -- 1990
         x"71",  x"f9",  x"a1",  x"80",  x"f3",  x"db",  x"89",  x"17", -- 1998
         x"0f",  x"d3",  x"89",  x"fb",  x"c9",  x"21",  x"a2",  x"b7", -- 19A0
         x"cb",  x"f6",  x"18",  x"e8",  x"0e",  x"20",  x"18",  x"d0", -- 19A8
         x"7f",  x"7f",  x"4c",  x"53",  x"54",  x"44",  x"45",  x"56", -- 19B0
         x"01",  x"cd",  x"8f",  x"fb",  x"cd",  x"a4",  x"c8",  x"c3", -- 19B8
         x"9c",  x"fb",  x"f5",  x"dd",  x"7e",  x"04",  x"f5",  x"dd", -- 19C0
         x"cb",  x"04",  x"ff",  x"d3",  x"86",  x"cd",  x"62",  x"ca", -- 19C8
         x"f1",  x"dd",  x"77",  x"04",  x"d3",  x"86",  x"f1",  x"c9", -- 19D0
         x"7f",  x"7f",  x"56",  x"32",  x"34",  x"44",  x"55",  x"50", -- 19D8
         x"01",  x"cd",  x"8f",  x"fb",  x"cd",  x"85",  x"c9",  x"dc", -- 19E0
         x"d1",  x"f4",  x"18",  x"d3",  x"cd",  x"8c",  x"e0",  x"dd", -- 19E8
         x"cb",  x"04",  x"7e",  x"20",  x"08",  x"e5",  x"21",  x"9c", -- 19F0
         x"fb",  x"e3",  x"cd",  x"8f",  x"fb",  x"c3",  x"12",  x"ca", -- 19F8
         x"c5",  x"f5",  x"0e",  x"05",  x"ed",  x"40",  x"cb",  x"50", -- 1A00
         x"20",  x"fa",  x"06",  x"01",  x"f3",  x"d3",  x"04",  x"18", -- 1A08
         x"0f",  x"c5",  x"f5",  x"0e",  x"90",  x"ed",  x"40",  x"cb", -- 1A10
         x"70",  x"20",  x"fa",  x"06",  x"80",  x"f3",  x"d3",  x"91", -- 1A18
         x"af",  x"ed",  x"79",  x"fb",  x"ed",  x"41",  x"f1",  x"c1", -- 1A20
         x"c9",  x"c5",  x"f5",  x"cd",  x"83",  x"fa",  x"c6",  x"0a", -- 1A28
         x"4f",  x"ed",  x"78",  x"e6",  x"04",  x"20",  x"03",  x"3c", -- 1A30
         x"18",  x"f7",  x"0d",  x"0d",  x"f1",  x"ed",  x"79",  x"c1", -- 1A38
         x"c9",  x"c5",  x"f5",  x"cd",  x"8b",  x"fa",  x"18",  x"e6", -- 1A40
         x"3e",  x"ee",  x"18",  x"03",  x"3a",  x"e8",  x"b7",  x"c5", -- 1A48
         x"d5",  x"57",  x"e6",  x"04",  x"0f",  x"0f",  x"c6",  x"0a", -- 1A50
         x"4f",  x"3e",  x"68",  x"a2",  x"5f",  x"ed",  x"78",  x"e6", -- 1A58
         x"01",  x"3e",  x"05",  x"f3",  x"ed",  x"79",  x"20",  x"0b", -- 1A60
         x"3e",  x"82",  x"b3",  x"ed",  x"79",  x"fb",  x"cd",  x"7c", -- 1A68
         x"e3",  x"30",  x"ea",  x"ed",  x"59",  x"fb",  x"38",  x"08", -- 1A70
         x"0d",  x"0d",  x"ed",  x"40",  x"3e",  x"7f",  x"b2",  x"a0", -- 1A78
         x"d1",  x"c1",  x"c9",  x"3a",  x"e1",  x"b7",  x"e6",  x"04", -- 1A80
         x"0f",  x"0f",  x"c9",  x"3a",  x"e8",  x"b7",  x"18",  x"f6", -- 1A88
         x"e5",  x"d5",  x"c5",  x"f5",  x"21",  x"00",  x"a8",  x"cd", -- 1A90
         x"86",  x"e3",  x"47",  x"0e",  x"80",  x"3e",  x"01",  x"ed", -- 1A98
         x"79",  x"d9",  x"d5",  x"c5",  x"db",  x"88",  x"47",  x"dd", -- 1AA0
         x"4e",  x"04",  x"dd",  x"cb",  x"04",  x"ff",  x"d3",  x"86", -- 1AA8
         x"d9",  x"21",  x"48",  x"d8",  x"f3",  x"db",  x"09",  x"cd", -- 1AB0
         x"4f",  x"f5",  x"cd",  x"b3",  x"e5",  x"fe",  x"0d",  x"28", -- 1AB8
         x"2d",  x"fe",  x"1b",  x"20",  x"0a",  x"cd",  x"48",  x"fa", -- 1AC0
         x"d6",  x"54",  x"28",  x"2e",  x"3d",  x"28",  x"74",  x"26", -- 1AC8
         x"b8",  x"68",  x"cd",  x"86",  x"e3",  x"21",  x"3b",  x"d8", -- 1AD0
         x"0e",  x"80",  x"f3",  x"cd",  x"4f",  x"f5",  x"ed",  x"79", -- 1AD8
         x"fb",  x"d9",  x"79",  x"dd",  x"77",  x"04",  x"d3",  x"86", -- 1AE0
         x"c1",  x"d1",  x"d9",  x"c3",  x"97",  x"e0",  x"f3",  x"dd", -- 1AE8
         x"36",  x"f2",  x"97",  x"dd",  x"36",  x"f3",  x"e3",  x"fb", -- 1AF0
         x"18",  x"d5",  x"21",  x"01",  x"b8",  x"cd",  x"86",  x"e3", -- 1AF8
         x"e6",  x"01",  x"07",  x"07",  x"d9",  x"57",  x"3e",  x"7b", -- 1B00
         x"a0",  x"b2",  x"57",  x"d9",  x"dd",  x"cb",  x"04",  x"bf", -- 1B08
         x"d3",  x"86",  x"cd",  x"48",  x"fa",  x"6f",  x"cd",  x"48", -- 1B10
         x"fa",  x"67",  x"cd",  x"48",  x"fa",  x"5f",  x"cd",  x"48", -- 1B18
         x"fa",  x"57",  x"cd",  x"48",  x"fa",  x"38",  x"14",  x"4f", -- 1B20
         x"d9",  x"7a",  x"d9",  x"f3",  x"d3",  x"88",  x"71",  x"d9", -- 1B28
         x"78",  x"d3",  x"88",  x"fb",  x"d9",  x"23",  x"1b",  x"7b", -- 1B30
         x"b2",  x"20",  x"e7",  x"dd",  x"cb",  x"04",  x"ff",  x"d3", -- 1B38
         x"86",  x"18",  x"8c",  x"cd",  x"48",  x"fa",  x"5f",  x"cd", -- 1B40
         x"48",  x"fa",  x"57",  x"21",  x"3b",  x"d8",  x"d9",  x"78", -- 1B48
         x"d9",  x"f6",  x"04",  x"f3",  x"cd",  x"4f",  x"f5",  x"d3", -- 1B50
         x"88",  x"dd",  x"cb",  x"04",  x"bf",  x"d3",  x"86",  x"ed", -- 1B58
         x"7b",  x"ae",  x"b7",  x"26",  x"b8",  x"68",  x"7e",  x"ed", -- 1B60
         x"79",  x"fb",  x"21",  x"69",  x"f2",  x"e5",  x"eb",  x"e9", -- 1B68
         x"cd",  x"9c",  x"fb",  x"f5",  x"3a",  x"01",  x"b8",  x"e6", -- 1B70
         x"01",  x"cc",  x"3f",  x"f0",  x"f1",  x"77",  x"18",  x"0c", -- 1B78
         x"cd",  x"9c",  x"fb",  x"3a",  x"01",  x"b8",  x"e6",  x"01", -- 1B80
         x"cc",  x"3f",  x"f0",  x"7e",  x"cd",  x"48",  x"f0",  x"f5", -- 1B88
         x"dd",  x"cb",  x"04",  x"ff",  x"18",  x"12",  x"cd",  x"8f", -- 1B90
         x"fb",  x"cd",  x"5c",  x"c1",  x"f5",  x"3a",  x"05",  x"b8", -- 1B98
         x"e6",  x"01",  x"20",  x"06",  x"dd",  x"cb",  x"04",  x"bf", -- 1BA0
         x"d3",  x"86",  x"f1",  x"c9",  x"cd",  x"8f",  x"fb",  x"cd", -- 1BA8
         x"db",  x"d2",  x"18",  x"e8",  x"7f",  x"7f",  x"44",  x"45", -- 1BB0
         x"56",  x"49",  x"43",  x"45",  x"01",  x"a7",  x"28",  x"15", -- 1BB8
         x"7d",  x"fe",  x"08",  x"d2",  x"d1",  x"f4",  x"cd",  x"d7", -- 1BC0
         x"fb",  x"da",  x"d1",  x"f4",  x"cd",  x"d2",  x"fb",  x"c3", -- 1BC8
         x"db",  x"f4",  x"3e",  x"fe",  x"21",  x"3e",  x"ff",  x"cd", -- 1BD0
         x"8f",  x"fb",  x"cd",  x"f2",  x"d5",  x"c3",  x"9c",  x"fb", -- 1BD8
         x"7f",  x"7f",  x"44",  x"49",  x"52",  x"20",  x"1f",  x"cd", -- 1BE0
         x"c9",  x"e4",  x"08",  x"c9",  x"7f",  x"7f",  x"43",  x"44", -- 1BE8
         x"20",  x"1f",  x"cd",  x"c9",  x"e4",  x"09",  x"c9",  x"7f", -- 1BF0
         x"7f",  x"45",  x"52",  x"41",  x"20",  x"1f",  x"cd",  x"c9", -- 1BF8
         x"e4",  x"0a",  x"c9",  x"7f",  x"7f",  x"52",  x"45",  x"4e", -- 1C00
         x"20",  x"1f",  x"cd",  x"c9",  x"e4",  x"0b",  x"c9",  x"57", -- 1C08
         x"77",  x"41",  x"61",  x"32",  x"22",  x"08",  x"19",  x"10", -- 1C10
         x"0c",  x"2d",  x"3d",  x"f2",  x"f8",  x"59",  x"79",  x"45", -- 1C18
         x"65",  x"53",  x"73",  x"33",  x"23",  x"5e",  x"5d",  x"01", -- 1C20
         x"0f",  x"3a",  x"2a",  x"f3",  x"f9",  x"58",  x"78",  x"54", -- 1C28
         x"74",  x"46",  x"66",  x"35",  x"25",  x"50",  x"70",  x"1f", -- 1C30
         x"02",  x"30",  x"40",  x"f5",  x"fb",  x"56",  x"76",  x"55", -- 1C38
         x"75",  x"48",  x"68",  x"37",  x"27",  x"4f",  x"6f",  x"1a", -- 1C40
         x"14",  x"39",  x"29",  x"03",  x"04",  x"4e",  x"6e",  x"49", -- 1C48
         x"69",  x"4a",  x"6a",  x"38",  x"28",  x"20",  x"5b",  x"4b", -- 1C50
         x"6b",  x"2c",  x"3c",  x"13",  x"1b",  x"4d",  x"6d",  x"5a", -- 1C58
         x"7a",  x"47",  x"67",  x"36",  x"26",  x"1c",  x"1d",  x"4c", -- 1C60
         x"6c",  x"2e",  x"3e",  x"f6",  x"fc",  x"42",  x"62",  x"52", -- 1C68
         x"72",  x"44",  x"64",  x"34",  x"24",  x"5f",  x"5c",  x"2b", -- 1C70
         x"3b",  x"2f",  x"3f",  x"f4",  x"fa",  x"43",  x"63",  x"51", -- 1C78
         x"71",  x"16",  x"05",  x"31",  x"21",  x"0a",  x"12",  x"0b", -- 1C80
         x"11",  x"09",  x"18",  x"f1",  x"f7",  x"0d",  x"0e",  x"bf", -- 1C88
         x"f4",  x"01",  x"e2",  x"78",  x"e2",  x"bf",  x"f4",  x"bf", -- 1C90
         x"f4",  x"ba",  x"e1",  x"bf",  x"f4",  x"8c",  x"e2",  x"e0", -- 1C98
         x"e1",  x"c9",  x"e1",  x"d2",  x"e1",  x"f0",  x"e1",  x"56", -- 1CA0
         x"e2",  x"66",  x"e2",  x"bf",  x"f4",  x"dc",  x"e1",  x"64", -- 1CA8
         x"e2",  x"f5",  x"e1",  x"fc",  x"e1",  x"bf",  x"f4",  x"d8", -- 1CB0
         x"e2",  x"bf",  x"f4",  x"bf",  x"f4",  x"bf",  x"f4",  x"ea", -- 1CB8
         x"e1",  x"66",  x"e2",  x"37",  x"e2",  x"51",  x"f9",  x"bf", -- 1CC0
         x"f4",  x"bf",  x"f4",  x"d0",  x"e1",  x"04",  x"e2",  x"c9", -- 1CC8
         x"4e",  x"4b",  x"45",  x"59",  x"24",  x"ca",  x"4f",  x"59", -- 1CD0
         x"53",  x"54",  x"d3",  x"54",  x"52",  x"49",  x"4e",  x"47", -- 1CD8
         x"24",  x"c9",  x"4e",  x"53",  x"54",  x"52",  x"d2",  x"45", -- 1CE0
         x"4e",  x"55",  x"4d",  x"42",  x"45",  x"52",  x"c4",  x"45", -- 1CE8
         x"4c",  x"45",  x"54",  x"45",  x"d0",  x"41",  x"55",  x"53", -- 1CF0
         x"45",  x"c2",  x"45",  x"45",  x"50",  x"d7",  x"49",  x"4e", -- 1CF8
         x"44",  x"4f",  x"57",  x"c2",  x"4f",  x"52",  x"44",  x"45", -- 1D00
         x"52",  x"c9",  x"4e",  x"4b",  x"d0",  x"41",  x"50",  x"45", -- 1D08
         x"52",  x"c1",  x"54",  x"c3",  x"4f",  x"4c",  x"4f",  x"52", -- 1D10
         x"d3",  x"4f",  x"55",  x"4e",  x"44",  x"d0",  x"53",  x"45", -- 1D18
         x"54",  x"d0",  x"52",  x"45",  x"53",  x"45",  x"54",  x"c2", -- 1D20
         x"4c",  x"4f",  x"41",  x"44",  x"d6",  x"50",  x"45",  x"45", -- 1D28
         x"4b",  x"d6",  x"50",  x"4f",  x"4b",  x"45",  x"cc",  x"4f", -- 1D30
         x"43",  x"41",  x"54",  x"45",  x"cb",  x"45",  x"59",  x"4c", -- 1D38
         x"49",  x"53",  x"54",  x"cb",  x"45",  x"59",  x"d3",  x"57", -- 1D40
         x"49",  x"54",  x"43",  x"48",  x"d0",  x"54",  x"45",  x"53", -- 1D48
         x"54",  x"c3",  x"4c",  x"4f",  x"53",  x"45",  x"cf",  x"50", -- 1D50
         x"45",  x"4e",  x"d2",  x"41",  x"4e",  x"44",  x"4f",  x"4d", -- 1D58
         x"49",  x"5a",  x"45",  x"d6",  x"47",  x"45",  x"54",  x"24", -- 1D60
         x"cc",  x"49",  x"4e",  x"45",  x"c3",  x"49",  x"52",  x"43", -- 1D68
         x"4c",  x"45",  x"c3",  x"53",  x"52",  x"4c",  x"49",  x"4e", -- 1D70
         x"c4",  x"45",  x"56",  x"49",  x"43",  x"45",  x"c6",  x"49", -- 1D78
         x"4c",  x"45",  x"53",  x"c3",  x"48",  x"44",  x"49",  x"52", -- 1D80
         x"80",  x"dd",  x"e9",  x"54",  x"ec",  x"43",  x"e6",  x"a5", -- 1D88
         x"ea",  x"a2",  x"e6",  x"81",  x"e8",  x"a5",  x"e8",  x"d5", -- 1D90
         x"e8",  x"f0",  x"e8",  x"21",  x"d4",  x"fb",  x"e9",  x"1c", -- 1D98
         x"ea",  x"48",  x"c3",  x"0d",  x"ea",  x"6b",  x"ea",  x"33", -- 1DA0
         x"ea",  x"30",  x"ea",  x"03",  x"ed",  x"48",  x"c3",  x"2f", -- 1DA8
         x"e9",  x"ac",  x"e9",  x"1a",  x"eb",  x"0f",  x"eb",  x"26", -- 1DB0
         x"eb",  x"48",  x"c3",  x"1c",  x"ec",  x"83",  x"ec",  x"7d", -- 1DB8
         x"ec",  x"48",  x"c3",  x"b8",  x"ec",  x"bd",  x"ec",  x"48", -- 1DC0
         x"c3",  x"e4",  x"ec",  x"29",  x"ed",  x"44",  x"ed",  x"ff", -- 1DC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1DD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1DD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1DE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1DE8
         x"16",  x"24",  x"37",  x"38",  x"06",  x"02",  x"07",  x"03", -- 1DF0
         x"80",  x"40",  x"20",  x"10",  x"08",  x"04",  x"02",  x"01", -- 1DF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"81",  x"ff", -- 1E00
         x"00",  x"00",  x"22",  x"72",  x"22",  x"3e",  x"00",  x"00", -- 1E08
         x"00",  x"32",  x"62",  x"fe",  x"62",  x"32",  x"00",  x"00", -- 1E10
         x"7e",  x"81",  x"b9",  x"a5",  x"b9",  x"a5",  x"b9",  x"81", -- 1E18
         x"55",  x"ff",  x"55",  x"ff",  x"55",  x"ff",  x"55",  x"ff", -- 1E20
         x"aa",  x"aa",  x"aa",  x"aa",  x"aa",  x"aa",  x"aa",  x"aa", -- 1E28
         x"ff",  x"00",  x"ff",  x"00",  x"ff",  x"00",  x"ff",  x"00", -- 1E30
         x"00",  x"00",  x"3c",  x"42",  x"42",  x"7e",  x"00",  x"00", -- 1E38
         x"00",  x"30",  x"60",  x"fe",  x"60",  x"30",  x"00",  x"00", -- 1E40
         x"00",  x"18",  x"0c",  x"fe",  x"0c",  x"18",  x"00",  x"00", -- 1E48
         x"10",  x"10",  x"10",  x"54",  x"7c",  x"38",  x"10",  x"00", -- 1E50
         x"10",  x"38",  x"7c",  x"54",  x"10",  x"10",  x"10",  x"00", -- 1E58
         x"70",  x"60",  x"50",  x"10",  x"10",  x"10",  x"7c",  x"00", -- 1E60
         x"00",  x"02",  x"12",  x"32",  x"7e",  x"30",  x"10",  x"00", -- 1E68
         x"aa",  x"55",  x"aa",  x"55",  x"aa",  x"55",  x"aa",  x"55", -- 1E70
         x"3e",  x"7c",  x"7c",  x"3e",  x"3e",  x"7c",  x"f8",  x"f8", -- 1E78
         x"38",  x"30",  x"28",  x"04",  x"04",  x"04",  x"04",  x"00", -- 1E80
         x"fe",  x"10",  x"38",  x"7c",  x"54",  x"10",  x"10",  x"00", -- 1E88
         x"10",  x"10",  x"54",  x"7c",  x"38",  x"10",  x"fe",  x"00", -- 1E90
         x"7e",  x"81",  x"9d",  x"a1",  x"99",  x"85",  x"b9",  x"81", -- 1E98
         x"00",  x"3c",  x"42",  x"5a",  x"5a",  x"42",  x"3c",  x"00", -- 1EA0
         x"88",  x"44",  x"22",  x"11",  x"88",  x"44",  x"22",  x"11", -- 1EA8
         x"00",  x"fe",  x"44",  x"e4",  x"4e",  x"44",  x"fe",  x"00", -- 1EB0
         x"11",  x"22",  x"44",  x"88",  x"11",  x"22",  x"44",  x"88", -- 1EB8
         x"02",  x"32",  x"1a",  x"fe",  x"1a",  x"32",  x"02",  x"00", -- 1EC0
         x"80",  x"98",  x"b0",  x"fe",  x"b0",  x"98",  x"80",  x"00", -- 1EC8
         x"00",  x"08",  x"7c",  x"06",  x"7c",  x"08",  x"00",  x"00", -- 1ED0
         x"cc",  x"cc",  x"33",  x"33",  x"cc",  x"cc",  x"33",  x"33", -- 1ED8
         x"7e",  x"81",  x"a1",  x"a1",  x"a1",  x"a1",  x"bd",  x"81", -- 1EE0
         x"7e",  x"81",  x"b9",  x"a5",  x"b9",  x"a5",  x"a5",  x"81", -- 1EE8
         x"7e",  x"81",  x"99",  x"a5",  x"a1",  x"a5",  x"99",  x"81", -- 1EF0
         x"00",  x"10",  x"3e",  x"60",  x"3e",  x"10",  x"00",  x"00", -- 1EF8
         x"3c",  x"42",  x"99",  x"a1",  x"a1",  x"99",  x"42",  x"3c", -- 1F00
         x"00",  x"00",  x"78",  x"0c",  x"7c",  x"cc",  x"76",  x"00", -- 1F08
         x"e0",  x"60",  x"7c",  x"66",  x"66",  x"66",  x"dc",  x"00", -- 1F10
         x"00",  x"00",  x"78",  x"cc",  x"c0",  x"cc",  x"78",  x"00", -- 1F18
         x"1c",  x"0c",  x"7c",  x"cc",  x"cc",  x"cc",  x"76",  x"00", -- 1F20
         x"00",  x"00",  x"78",  x"cc",  x"fc",  x"c0",  x"78",  x"00", -- 1F28
         x"38",  x"6c",  x"60",  x"f0",  x"60",  x"60",  x"f0",  x"00", -- 1F30
         x"00",  x"00",  x"76",  x"cc",  x"cc",  x"7c",  x"0c",  x"f8", -- 1F38
         x"e0",  x"60",  x"6c",  x"76",  x"66",  x"66",  x"e6",  x"00", -- 1F40
         x"30",  x"00",  x"70",  x"30",  x"30",  x"30",  x"fc",  x"00", -- 1F48
         x"0c",  x"00",  x"1c",  x"0c",  x"0c",  x"cc",  x"cc",  x"78", -- 1F50
         x"e0",  x"60",  x"66",  x"6c",  x"78",  x"6c",  x"e6",  x"00", -- 1F58
         x"70",  x"30",  x"30",  x"30",  x"30",  x"30",  x"fc",  x"00", -- 1F60
         x"00",  x"00",  x"cc",  x"fe",  x"fe",  x"d6",  x"c6",  x"00", -- 1F68
         x"00",  x"00",  x"f8",  x"cc",  x"cc",  x"cc",  x"cc",  x"00", -- 1F70
         x"00",  x"00",  x"78",  x"cc",  x"cc",  x"cc",  x"78",  x"00", -- 1F78
         x"00",  x"00",  x"dc",  x"66",  x"66",  x"7c",  x"60",  x"f0", -- 1F80
         x"00",  x"00",  x"76",  x"cc",  x"cc",  x"7c",  x"0c",  x"1e", -- 1F88
         x"00",  x"00",  x"dc",  x"76",  x"66",  x"60",  x"f0",  x"00", -- 1F90
         x"00",  x"00",  x"7c",  x"c0",  x"78",  x"0c",  x"f8",  x"00", -- 1F98
         x"10",  x"30",  x"7c",  x"30",  x"30",  x"34",  x"18",  x"00", -- 1FA0
         x"00",  x"00",  x"cc",  x"cc",  x"cc",  x"cc",  x"76",  x"00", -- 1FA8
         x"00",  x"00",  x"cc",  x"cc",  x"cc",  x"78",  x"30",  x"00", -- 1FB0
         x"00",  x"00",  x"c6",  x"d6",  x"fe",  x"fe",  x"6c",  x"00", -- 1FB8
         x"00",  x"00",  x"c6",  x"6c",  x"38",  x"6c",  x"c6",  x"00", -- 1FC0
         x"00",  x"00",  x"cc",  x"cc",  x"cc",  x"7c",  x"0c",  x"f8", -- 1FC8
         x"00",  x"00",  x"fc",  x"98",  x"30",  x"64",  x"fc",  x"00", -- 1FD0
         x"6c",  x"00",  x"78",  x"0c",  x"7c",  x"cc",  x"76",  x"00", -- 1FD8
         x"cc",  x"00",  x"78",  x"cc",  x"cc",  x"cc",  x"78",  x"00", -- 1FE0
         x"cc",  x"00",  x"cc",  x"cc",  x"cc",  x"cc",  x"76",  x"00", -- 1FE8
         x"3c",  x"66",  x"66",  x"6c",  x"66",  x"66",  x"6c",  x"f0", -- 1FF0
         x"ff",  x"81",  x"81",  x"81",  x"81",  x"81",  x"81",  x"ff"  -- 1FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
