library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity user47_c is
    generic(
        ADDR_WIDTH   : integer := 15
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end user47_c;

architecture rtl of user47_c is
    type rom32768x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom32768x8 := (
         x"00",  x"00",  x"00",  x"00",  x"00",  x"22",  x"22",  x"22", -- 0000
         x"22",  x"22",  x"00",  x"ff",  x"ec",  x"80",  x"00",  x"00", -- 0008
         x"ff",  x"73",  x"10",  x"00",  x"07",  x"65",  x"11",  x"11", -- 0010
         x"00",  x"00",  x"01",  x"e6",  x"20",  x"00",  x"00",  x"f0", -- 0018
         x"20",  x"20",  x"00",  x"88",  x"f0",  x"00",  x"00",  x"00", -- 0020
         x"00",  x"26",  x"f6",  x"20",  x"00",  x"00",  x"46",  x"f6", -- 0028
         x"40",  x"00",  x"02",  x"22",  x"22",  x"72",  x"00",  x"02", -- 0030
         x"72",  x"22",  x"22",  x"00",  x"0e",  x"ca",  x"22",  x"27", -- 0038
         x"00",  x"01",  x"11",  x"5f",  x"40",  x"00",  x"01",  x"11", -- 0040
         x"13",  x"73",  x"00",  x"01",  x"24",  x"a5",  x"24",  x"80", -- 0048
         x"07",  x"55",  x"57",  x"00",  x"00",  x"01",  x"31",  x"11", -- 0050
         x"00",  x"00",  x"07",  x"17",  x"47",  x"00",  x"00",  x"07", -- 0058
         x"17",  x"17",  x"00",  x"00",  x"04",  x"57",  x"11",  x"00", -- 0060
         x"00",  x"07",  x"47",  x"17",  x"00",  x"00",  x"07",  x"47", -- 0068
         x"57",  x"00",  x"00",  x"07",  x"11",  x"11",  x"00",  x"00", -- 0070
         x"07",  x"57",  x"57",  x"00",  x"00",  x"07",  x"57",  x"17", -- 0078
         x"00",  x"00",  x"0f",  x"f0",  x"ff",  x"0f",  x"f0",  x"96", -- 0080
         x"69",  x"96",  x"69",  x"00",  x"00",  x"13",  x"73",  x"10", -- 0088
         x"00",  x"02",  x"72",  x"22",  x"20",  x"00",  x"00",  x"46", -- 0090
         x"76",  x"40",  x"00",  x"02",  x"22",  x"27",  x"20",  x"00", -- 0098
         x"00",  x"00",  x"00",  x"00",  x"00",  x"02",  x"77",  x"22", -- 00A0
         x"02",  x"00",  x"05",  x"50",  x"00",  x"00",  x"00",  x"00", -- 00A8
         x"57",  x"57",  x"50",  x"00",  x"02",  x"76",  x"23",  x"72", -- 00B0
         x"00",  x"00",  x"51",  x"22",  x"45",  x"00",  x"00",  x"25", -- 00B8
         x"25",  x"43",  x"00",  x"02",  x"20",  x"00",  x"00",  x"00", -- 00C0
         x"01",  x"22",  x"22",  x"21",  x"00",  x"04",  x"22",  x"22", -- 00C8
         x"24",  x"00",  x"00",  x"05",  x"25",  x"00",  x"00",  x"00", -- 00D0
         x"02",  x"72",  x"00",  x"00",  x"00",  x"00",  x"00",  x"22", -- 00D8
         x"40",  x"00",  x"00",  x"70",  x"00",  x"00",  x"00",  x"00", -- 00E0
         x"00",  x"02",  x"00",  x"01",  x"12",  x"22",  x"44",  x"00", -- 00E8
         x"02",  x"55",  x"55",  x"52",  x"00",  x"01",  x"35",  x"11", -- 00F0
         x"11",  x"00",  x"02",  x"55",  x"12",  x"47",  x"00",  x"02", -- 00F8
         x"51",  x"21",  x"52",  x"00",  x"04",  x"55",  x"71",  x"11", -- 0100
         x"00",  x"07",  x"44",  x"71",  x"52",  x"00",  x"02",  x"44", -- 0108
         x"65",  x"52",  x"00",  x"07",  x"11",  x"12",  x"22",  x"00", -- 0110
         x"02",  x"55",  x"25",  x"52",  x"00",  x"02",  x"55",  x"31", -- 0118
         x"52",  x"00",  x"00",  x"02",  x"00",  x"20",  x"00",  x"00", -- 0120
         x"02",  x"00",  x"22",  x"40",  x"00",  x"12",  x"42",  x"10", -- 0128
         x"00",  x"00",  x"07",  x"07",  x"00",  x"00",  x"00",  x"42", -- 0130
         x"12",  x"40",  x"00",  x"02",  x"51",  x"22",  x"02",  x"00", -- 0138
         x"06",  x"51",  x"25",  x"53",  x"00",  x"02",  x"55",  x"75", -- 0140
         x"55",  x"00",  x"06",  x"55",  x"65",  x"56",  x"00",  x"02", -- 0148
         x"54",  x"44",  x"52",  x"00",  x"06",  x"55",  x"55",  x"56", -- 0150
         x"00",  x"07",  x"44",  x"64",  x"47",  x"00",  x"07",  x"44", -- 0158
         x"64",  x"44",  x"00",  x"02",  x"54",  x"45",  x"53",  x"00", -- 0160
         x"05",  x"55",  x"75",  x"55",  x"00",  x"07",  x"22",  x"22", -- 0168
         x"27",  x"00",  x"07",  x"11",  x"11",  x"52",  x"00",  x"05", -- 0170
         x"56",  x"46",  x"55",  x"00",  x"04",  x"44",  x"44",  x"47", -- 0178
         x"00",  x"05",  x"77",  x"55",  x"55",  x"00",  x"06",  x"55", -- 0180
         x"55",  x"55",  x"00",  x"07",  x"55",  x"55",  x"57",  x"00", -- 0188
         x"06",  x"55",  x"64",  x"44",  x"00",  x"07",  x"55",  x"55", -- 0190
         x"77",  x"10",  x"06",  x"55",  x"65",  x"55",  x"00",  x"02", -- 0198
         x"54",  x"21",  x"52",  x"00",  x"07",  x"22",  x"22",  x"22", -- 01A0
         x"00",  x"05",  x"55",  x"55",  x"57",  x"00",  x"05",  x"55", -- 01A8
         x"55",  x"52",  x"00",  x"05",  x"55",  x"57",  x"75",  x"00", -- 01B0
         x"05",  x"55",  x"25",  x"55",  x"00",  x"05",  x"55",  x"72", -- 01B8
         x"22",  x"00",  x"07",  x"11",  x"24",  x"47",  x"00",  x"07", -- 01C0
         x"44",  x"44",  x"47",  x"00",  x"04",  x"42",  x"22",  x"11", -- 01C8
         x"00",  x"07",  x"11",  x"11",  x"17",  x"00",  x"00",  x"25", -- 01D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"70", -- 01D8
         x"00",  x"21",  x"00",  x"00",  x"00",  x"00",  x"02",  x"55", -- 01E0
         x"53",  x"00",  x"04",  x"46",  x"55",  x"56",  x"00",  x"00", -- 01E8
         x"03",  x"44",  x"43",  x"00",  x"01",  x"13",  x"55",  x"53", -- 01F0
         x"00",  x"00",  x"02",  x"57",  x"47",  x"00",  x"02",  x"54", -- 01F8
         x"64",  x"44",  x"40",  x"00",  x"03",  x"55",  x"31",  x"60", -- 0200
         x"04",  x"46",  x"55",  x"55",  x"00",  x"00",  x"20",  x"22", -- 0208
         x"22",  x"00",  x"00",  x"20",  x"22",  x"22",  x"60",  x"04", -- 0210
         x"45",  x"56",  x"55",  x"00",  x"04",  x"44",  x"44",  x"52", -- 0218
         x"00",  x"00",  x"05",  x"75",  x"55",  x"00",  x"00",  x"02", -- 0220
         x"55",  x"55",  x"00",  x"00",  x"02",  x"55",  x"52",  x"00", -- 0228
         x"00",  x"02",  x"55",  x"64",  x"40",  x"00",  x"02",  x"55", -- 0230
         x"31",  x"10",  x"00",  x"06",  x"54",  x"44",  x"00",  x"00", -- 0238
         x"03",  x"42",  x"16",  x"00",  x"02",  x"27",  x"22",  x"21", -- 0240
         x"00",  x"00",  x"05",  x"55",  x"57",  x"00",  x"00",  x"05", -- 0248
         x"55",  x"52",  x"00",  x"00",  x"05",  x"57",  x"75",  x"00", -- 0250
         x"00",  x"05",  x"52",  x"55",  x"00",  x"00",  x"05",  x"55", -- 0258
         x"31",  x"60",  x"00",  x"07",  x"12",  x"47",  x"00",  x"03", -- 0260
         x"22",  x"42",  x"23",  x"00",  x"02",  x"22",  x"22",  x"22", -- 0268
         x"00",  x"06",  x"22",  x"12",  x"26",  x"00",  x"07",  x"00", -- 0270
         x"00",  x"00",  x"00",  x"07",  x"77",  x"77",  x"77",  x"70", -- 0278
         x"02",  x"54",  x"44",  x"52",  x"40",  x"00",  x"50",  x"55", -- 0280
         x"57",  x"00",  x"12",  x"02",  x"57",  x"43",  x"00",  x"02", -- 0288
         x"50",  x"25",  x"53",  x"00",  x"00",  x"50",  x"25",  x"53", -- 0290
         x"00",  x"04",  x"20",  x"25",  x"53",  x"00",  x"00",  x"20", -- 0298
         x"25",  x"53",  x"00",  x"00",  x"03",  x"44",  x"43",  x"40", -- 02A0
         x"25",  x"02",  x"57",  x"47",  x"00",  x"05",  x"02",  x"57", -- 02A8
         x"47",  x"00",  x"42",  x"02",  x"57",  x"47",  x"00",  x"05", -- 02B0
         x"02",  x"22",  x"22",  x"00",  x"25",  x"02",  x"22",  x"22", -- 02B8
         x"00",  x"04",  x"20",  x"22",  x"22",  x"00",  x"05",  x"25", -- 02C0
         x"57",  x"55",  x"00",  x"25",  x"25",  x"57",  x"55",  x"00", -- 02C8
         x"12",  x"07",  x"46",  x"47",  x"00",  x"00",  x"05",  x"37", -- 02D0
         x"65",  x"00",  x"07",  x"aa",  x"fa",  x"ab",  x"00",  x"02", -- 02D8
         x"50",  x"25",  x"52",  x"00",  x"00",  x"50",  x"25",  x"52", -- 02E0
         x"00",  x"04",  x"20",  x"25",  x"52",  x"00",  x"02",  x"50", -- 02E8
         x"55",  x"53",  x"00",  x"04",  x"20",  x"55",  x"53",  x"00", -- 02F0
         x"05",  x"05",  x"55",  x"31",  x"60",  x"05",  x"07",  x"55", -- 02F8
         x"57",  x"00",  x"05",  x"05",  x"55",  x"57",  x"00",  x"00", -- 0300
         x"27",  x"66",  x"67",  x"20",  x"02",  x"54",  x"64",  x"47", -- 0308
         x"00",  x"05",  x"52",  x"72",  x"72",  x"00",  x"0c",  x"ac", -- 0310
         x"ab",  x"ab",  x"00",  x"00",  x"32",  x"72",  x"22",  x"60", -- 0318
         x"01",  x"20",  x"25",  x"53",  x"00",  x"01",  x"20",  x"22", -- 0320
         x"22",  x"00",  x"01",  x"20",  x"25",  x"52",  x"00",  x"01", -- 0328
         x"20",  x"55",  x"57",  x"00",  x"00",  x"70",  x"25",  x"55", -- 0330
         x"00",  x"07",  x"06",  x"55",  x"55",  x"00",  x"00",  x"25", -- 0338
         x"55",  x"30",  x"70",  x"00",  x"25",  x"55",  x"20",  x"70", -- 0340
         x"02",  x"02",  x"24",  x"52",  x"00",  x"00",  x"f8",  x"00", -- 0348
         x"00",  x"00",  x"00",  x"f1",  x"00",  x"00",  x"00",  x"44", -- 0350
         x"52",  x"51",  x"27",  x"00",  x"44",  x"41",  x"25",  x"71", -- 0358
         x"00",  x"02",  x"02",  x"27",  x"72",  x"00",  x"00",  x"05", -- 0360
         x"a5",  x"00",  x"00",  x"00",  x"0a",  x"5a",  x"00",  x"00", -- 0368
         x"05",  x"05",  x"05",  x"05",  x"05",  x"aa",  x"55",  x"aa", -- 0370
         x"55",  x"aa",  x"a5",  x"a5",  x"a5",  x"a5",  x"a5",  x"22", -- 0378
         x"22",  x"22",  x"22",  x"22",  x"22",  x"2e",  x"22",  x"22", -- 0380
         x"22",  x"22",  x"e2",  x"e2",  x"22",  x"22",  x"66",  x"6e", -- 0388
         x"66",  x"66",  x"66",  x"00",  x"0e",  x"66",  x"66",  x"66", -- 0390
         x"00",  x"e2",  x"e2",  x"22",  x"22",  x"66",  x"e2",  x"e6", -- 0398
         x"66",  x"66",  x"66",  x"66",  x"66",  x"66",  x"66",  x"00", -- 03A0
         x"e2",  x"e6",  x"66",  x"66",  x"66",  x"e2",  x"e0",  x"00", -- 03A8
         x"00",  x"66",  x"6e",  x"00",  x"00",  x"00",  x"22",  x"e2", -- 03B0
         x"e0",  x"00",  x"00",  x"00",  x"0e",  x"22",  x"22",  x"22", -- 03B8
         x"22",  x"23",  x"00",  x"00",  x"00",  x"22",  x"2f",  x"00", -- 03C0
         x"00",  x"00",  x"00",  x"0f",  x"22",  x"22",  x"22",  x"22", -- 03C8
         x"23",  x"22",  x"22",  x"22",  x"00",  x"0f",  x"00",  x"00", -- 03D0
         x"00",  x"22",  x"2f",  x"22",  x"22",  x"22",  x"22",  x"32", -- 03D8
         x"32",  x"22",  x"22",  x"66",  x"67",  x"66",  x"66",  x"66", -- 03E0
         x"66",  x"74",  x"70",  x"00",  x"00",  x"00",  x"74",  x"76", -- 03E8
         x"66",  x"66",  x"66",  x"f0",  x"f0",  x"00",  x"00",  x"00", -- 03F0
         x"f0",  x"f6",  x"66",  x"66",  x"66",  x"74",  x"76",  x"66", -- 03F8
         x"66",  x"00",  x"f0",  x"f0",  x"00",  x"00",  x"66",  x"f0", -- 0400
         x"f6",  x"66",  x"66",  x"22",  x"f0",  x"f0",  x"00",  x"00", -- 0408
         x"66",  x"6f",  x"00",  x"00",  x"00",  x"00",  x"f0",  x"f2", -- 0410
         x"22",  x"22",  x"00",  x"0f",  x"66",  x"66",  x"66",  x"66", -- 0418
         x"67",  x"00",  x"00",  x"00",  x"22",  x"32",  x"30",  x"00", -- 0420
         x"00",  x"00",  x"32",  x"32",  x"22",  x"22",  x"00",  x"07", -- 0428
         x"66",  x"66",  x"66",  x"66",  x"6f",  x"66",  x"66",  x"66", -- 0430
         x"22",  x"f2",  x"f2",  x"22",  x"22",  x"22",  x"2e",  x"00", -- 0438
         x"00",  x"00",  x"00",  x"03",  x"22",  x"22",  x"22",  x"ff", -- 0440
         x"ff",  x"ff",  x"ff",  x"ff",  x"00",  x"00",  x"0f",  x"ff", -- 0448
         x"ff",  x"cc",  x"cc",  x"cc",  x"cc",  x"cc",  x"33",  x"33", -- 0450
         x"33",  x"33",  x"33",  x"ff",  x"ff",  x"f0",  x"00",  x"00", -- 0458
         x"00",  x"00",  x"16",  x"61",  x"00",  x"02",  x"55",  x"65", -- 0460
         x"56",  x"40",  x"07",  x"55",  x"44",  x"44",  x"00",  x"00", -- 0468
         x"00",  x"75",  x"55",  x"00",  x"07",  x"42",  x"12",  x"47", -- 0470
         x"00",  x"00",  x"01",  x"25",  x"52",  x"00",  x"00",  x"05", -- 0478
         x"55",  x"57",  x"44",  x"00",  x"07",  x"22",  x"24",  x"00", -- 0480
         x"07",  x"25",  x"55",  x"27",  x"00",  x"02",  x"55",  x"75", -- 0488
         x"52",  x"00",  x"02",  x"55",  x"52",  x"25",  x"00",  x"00", -- 0490
         x"34",  x"25",  x"52",  x"00",  x"00",  x"00",  x"6f",  x"60", -- 0498
         x"00",  x"07",  x"55",  x"75",  x"57",  x"00",  x"00",  x"34", -- 04A0
         x"74",  x"30",  x"00",  x"00",  x"25",  x"55",  x"55",  x"00", -- 04A8
         x"00",  x"70",  x"70",  x"70",  x"00",  x"00",  x"27",  x"20", -- 04B0
         x"07",  x"00",  x"04",  x"21",  x"24",  x"07",  x"00",  x"01", -- 04B8
         x"24",  x"21",  x"07",  x"00",  x"02",  x"54",  x"44",  x"42", -- 04C0
         x"22",  x"22",  x"11",  x"11",  x"52",  x"00",  x"00",  x"20", -- 04C8
         x"70",  x"20",  x"00",  x"00",  x"63",  x"06",  x"30",  x"00", -- 04D0
         x"02",  x"52",  x"00",  x"00",  x"00",  x"00",  x"02",  x"20", -- 04D8
         x"00",  x"00",  x"00",  x"00",  x"20",  x"00",  x"00",  x"03", -- 04E0
         x"22",  x"e6",  x"44",  x"00",  x"06",  x"55",  x"00",  x"00", -- 04E8
         x"00",  x"02",  x"51",  x"27",  x"00",  x"00",  x"00",  x"00", -- 04F0
         x"33",  x"00",  x"00",  x"0f",  x"99",  x"99",  x"99",  x"f0", -- 04F8
         x"03",  x"42",  x"52",  x"16",  x"00",  x"05",  x"25",  x"57", -- 0500
         x"55",  x"00",  x"05",  x"07",  x"55",  x"57",  x"00",  x"05", -- 0508
         x"05",  x"55",  x"57",  x"00",  x"00",  x"21",  x"00",  x"00", -- 0510
         x"00",  x"00",  x"50",  x"25",  x"53",  x"00",  x"00",  x"50", -- 0518
         x"25",  x"52",  x"00",  x"00",  x"50",  x"55",  x"57",  x"00", -- 0520
         x"02",  x"55",  x"65",  x"56",  x"40",  x"06",  x"51",  x"25", -- 0528
         x"53",  x"00",  x"0f",  x"ff",  x"ff",  x"ff",  x"f0",  x"02", -- 0530
         x"22",  x"22",  x"22",  x"00",  x"00",  x"f1",  x"00",  x"00", -- 0538
         x"00",  x"06",  x"9f",  x"df",  x"96",  x"00",  x"00",  x"50", -- 0540
         x"25",  x"53",  x"00",  x"00",  x"50",  x"25",  x"52",  x"00", -- 0548
         x"00",  x"50",  x"55",  x"57",  x"00",  x"02",  x"55",  x"65", -- 0550
         x"56",  x"40",  x"cd",  x"ea",  x"ca",  x"c3",  x"9c",  x"cb", -- 0558
         x"f5",  x"cd",  x"03",  x"f0",  x"33",  x"38",  x"1f",  x"d5", -- 0560
         x"3a",  x"9c",  x"b7",  x"83",  x"5f",  x"d5",  x"3a",  x"9d", -- 0568
         x"b7",  x"82",  x"87",  x"87",  x"87",  x"6f",  x"26",  x"00", -- 0570
         x"29",  x"54",  x"5d",  x"29",  x"29",  x"19",  x"d1",  x"16", -- 0578
         x"ad",  x"19",  x"d1",  x"f1",  x"a7",  x"c9",  x"f1",  x"37", -- 0580
         x"c9",  x"d5",  x"ed",  x"5b",  x"9c",  x"b7",  x"19",  x"d1", -- 0588
         x"cb",  x"3d",  x"f5",  x"3e",  x"80",  x"85",  x"44",  x"67", -- 0590
         x"78",  x"87",  x"87",  x"87",  x"80",  x"80",  x"c6",  x"06", -- 0598
         x"6f",  x"f1",  x"c9",  x"e5",  x"21",  x"a2",  x"b7",  x"cb", -- 05A0
         x"de",  x"cd",  x"36",  x"c6",  x"cb",  x"9e",  x"e1",  x"c9", -- 05A8
         x"af",  x"be",  x"c8",  x"77",  x"e5",  x"d5",  x"c5",  x"f5", -- 05B0
         x"21",  x"3e",  x"00",  x"cb",  x"6e",  x"20",  x"09",  x"cb", -- 05B8
         x"76",  x"28",  x"36",  x"21",  x"2d",  x"c5",  x"18",  x"03", -- 05C0
         x"21",  x"00",  x"c5",  x"fe",  x"40",  x"28",  x"36",  x"01", -- 05C8
         x"05",  x"00",  x"fe",  x"5b",  x"28",  x"2e",  x"09",  x"fe", -- 05D0
         x"5c",  x"28",  x"29",  x"09",  x"fe",  x"5d",  x"28",  x"24", -- 05D8
         x"09",  x"fe",  x"60",  x"28",  x"1f",  x"09",  x"fe",  x"7b", -- 05E0
         x"28",  x"1a",  x"09",  x"fe",  x"7c",  x"28",  x"15",  x"09", -- 05E8
         x"fe",  x"7d",  x"28",  x"10",  x"09",  x"fe",  x"7e",  x"28", -- 05F0
         x"0b",  x"26",  x"00",  x"6f",  x"44",  x"4f",  x"29",  x"29", -- 05F8
         x"09",  x"01",  x"00",  x"c0",  x"09",  x"eb",  x"cd",  x"89", -- 0600
         x"c5",  x"06",  x"05",  x"c5",  x"f5",  x"1a",  x"13",  x"47", -- 0608
         x"07",  x"07",  x"07",  x"07",  x"4f",  x"f1",  x"38",  x"0d", -- 0610
         x"ed",  x"6f",  x"79",  x"ed",  x"67",  x"23",  x"ed",  x"6f", -- 0618
         x"78",  x"ed",  x"67",  x"18",  x"0b",  x"ed",  x"67",  x"79", -- 0620
         x"ed",  x"6f",  x"23",  x"ed",  x"67",  x"78",  x"ed",  x"6f", -- 0628
         x"23",  x"c1",  x"10",  x"d7",  x"18",  x"36",  x"e5",  x"d5", -- 0630
         x"c5",  x"f5",  x"cd",  x"71",  x"c6",  x"ed",  x"53",  x"a0", -- 0638
         x"b7",  x"18",  x"29",  x"e5",  x"d5",  x"c5",  x"f5",  x"ed", -- 0640
         x"5b",  x"a0",  x"b7",  x"cd",  x"60",  x"c5",  x"7e",  x"a7", -- 0648
         x"f5",  x"eb",  x"cd",  x"89",  x"c5",  x"06",  x"0a",  x"0e", -- 0650
         x"f0",  x"30",  x"02",  x"0e",  x"0f",  x"f1",  x"20",  x"06", -- 0658
         x"3e",  x"08",  x"85",  x"6f",  x"06",  x"02",  x"7e",  x"a9", -- 0660
         x"77",  x"23",  x"10",  x"fa",  x"f1",  x"c1",  x"d1",  x"e1", -- 0668
         x"c9",  x"ed",  x"5b",  x"a0",  x"b7",  x"fe",  x"20",  x"30", -- 0670
         x"14",  x"21",  x"a2",  x"b7",  x"cb",  x"5e",  x"20",  x"0d", -- 0678
         x"87",  x"21",  x"14",  x"df",  x"4f",  x"06",  x"00",  x"09", -- 0680
         x"7e",  x"23",  x"66",  x"6f",  x"e9",  x"cd",  x"60",  x"c5", -- 0688
         x"d8",  x"77",  x"cd",  x"b4",  x"c5",  x"3a",  x"9e",  x"b7", -- 0690
         x"3d",  x"bb",  x"28",  x"03",  x"1c",  x"18",  x"0f",  x"3a", -- 0698
         x"9f",  x"b7",  x"3d",  x"ba",  x"20",  x"05",  x"cd",  x"f6", -- 06A0
         x"c6",  x"d8",  x"3e",  x"14",  x"1e",  x"00",  x"7b",  x"e6", -- 06A8
         x"07",  x"c8",  x"cd",  x"60",  x"c5",  x"7e",  x"b7",  x"c0", -- 06B0
         x"2b",  x"7e",  x"b7",  x"28",  x"d8",  x"c9",  x"cd",  x"95", -- 06B8
         x"c6",  x"d8",  x"cd",  x"60",  x"c5",  x"7e",  x"fe",  x"21", -- 06C0
         x"30",  x"f4",  x"cd",  x"60",  x"c5",  x"7e",  x"fe",  x"21", -- 06C8
         x"d0",  x"cd",  x"95",  x"c6",  x"d8",  x"18",  x"f3",  x"3a", -- 06D0
         x"9f",  x"b7",  x"3d",  x"ba",  x"20",  x"05",  x"cd",  x"f6", -- 06D8
         x"c6",  x"d8",  x"3e",  x"14",  x"cd",  x"60",  x"c5",  x"7e", -- 06E0
         x"fe",  x"20",  x"d0",  x"7b",  x"a7",  x"c8",  x"2b",  x"7e", -- 06E8
         x"fe",  x"20",  x"d0",  x"1d",  x"18",  x"f5",  x"d5",  x"2a", -- 06F0
         x"1a",  x"00",  x"ed",  x"5b",  x"1e",  x"00",  x"a7",  x"ed", -- 06F8
         x"52",  x"d1",  x"37",  x"c8",  x"d5",  x"11",  x"00",  x"00", -- 0700
         x"cd",  x"60",  x"c5",  x"cd",  x"2b",  x"d7",  x"38",  x"24", -- 0708
         x"cd",  x"a4",  x"c7",  x"ed",  x"5b",  x"9e",  x"b7",  x"15", -- 0710
         x"1e",  x"00",  x"cd",  x"60",  x"c5",  x"ed",  x"4b",  x"1e", -- 0718
         x"00",  x"e5",  x"2a",  x"1a",  x"00",  x"a7",  x"ed",  x"42", -- 0720
         x"e1",  x"c4",  x"88",  x"d7",  x"2a",  x"12",  x"00",  x"23", -- 0728
         x"22",  x"12",  x"00",  x"a7",  x"d1",  x"c9",  x"7a",  x"a7", -- 0730
         x"20",  x"05",  x"cd",  x"42",  x"c7",  x"d8",  x"3e",  x"15", -- 0738
         x"18",  x"a2",  x"d5",  x"2a",  x"1c",  x"00",  x"ed",  x"5b", -- 0740
         x"18",  x"00",  x"a7",  x"ed",  x"52",  x"d1",  x"37",  x"c8", -- 0748
         x"d5",  x"2a",  x"1c",  x"00",  x"e5",  x"ed",  x"5b",  x"9e", -- 0750
         x"b7",  x"15",  x"1e",  x"00",  x"cd",  x"60",  x"c5",  x"cd", -- 0758
         x"2b",  x"d7",  x"d1",  x"d4",  x"e8",  x"d6",  x"d1",  x"d5", -- 0760
         x"cd",  x"fe",  x"c7",  x"2a",  x"1c",  x"00",  x"06",  x"02", -- 0768
         x"2b",  x"cd",  x"86",  x"00",  x"fe",  x"0d",  x"20",  x"f8", -- 0770
         x"10",  x"f6",  x"23",  x"cd",  x"86",  x"00",  x"fe",  x"0a", -- 0778
         x"28",  x"f8",  x"22",  x"1c",  x"00",  x"2a",  x"1e",  x"00", -- 0780
         x"e5",  x"11",  x"00",  x"00",  x"cd",  x"60",  x"c5",  x"ed", -- 0788
         x"4b",  x"1c",  x"00",  x"cd",  x"88",  x"d7",  x"e1",  x"22", -- 0790
         x"1e",  x"00",  x"2a",  x"12",  x"00",  x"2b",  x"22",  x"12", -- 0798
         x"00",  x"d1",  x"a7",  x"c9",  x"06",  x"16",  x"3e",  x"16", -- 07A0
         x"90",  x"d8",  x"67",  x"2e",  x"00",  x"78",  x"87",  x"4f", -- 07A8
         x"87",  x"87",  x"81",  x"4f",  x"c5",  x"cd",  x"89",  x"c5", -- 07B0
         x"54",  x"5d",  x"7d",  x"c6",  x"0a",  x"6f",  x"3e",  x"28", -- 07B8
         x"e5",  x"d5",  x"c5",  x"06",  x"00",  x"ed",  x"b0",  x"eb", -- 07C0
         x"06",  x"0a",  x"36",  x"00",  x"23",  x"10",  x"fb",  x"c1", -- 07C8
         x"d1",  x"e1",  x"14",  x"24",  x"3d",  x"20",  x"e9",  x"c1", -- 07D0
         x"06",  x"00",  x"cb",  x"21",  x"cb",  x"10",  x"cb",  x"21", -- 07D8
         x"cb",  x"10",  x"cb",  x"21",  x"cb",  x"10",  x"21",  x"80", -- 07E0
         x"b4",  x"ed",  x"42",  x"54",  x"5d",  x"c5",  x"01",  x"50", -- 07E8
         x"00",  x"09",  x"c1",  x"ed",  x"b0",  x"eb",  x"06",  x"50", -- 07F0
         x"af",  x"77",  x"23",  x"10",  x"fc",  x"c9",  x"06",  x"16", -- 07F8
         x"3e",  x"16",  x"90",  x"d8",  x"78",  x"87",  x"4f",  x"87", -- 0800
         x"87",  x"81",  x"4f",  x"06",  x"00",  x"16",  x"80",  x"62", -- 0808
         x"3e",  x"28",  x"1e",  x"ff",  x"2e",  x"f5",  x"c5",  x"0c", -- 0810
         x"0d",  x"28",  x"02",  x"ed",  x"b8",  x"06",  x"0a",  x"23", -- 0818
         x"36",  x"00",  x"10",  x"fb",  x"c1",  x"14",  x"24",  x"3d", -- 0820
         x"20",  x"e8",  x"11",  x"cf",  x"b4",  x"21",  x"7f",  x"b4", -- 0828
         x"0c",  x"0d",  x"28",  x"0e",  x"cb",  x"21",  x"cb",  x"10", -- 0830
         x"cb",  x"21",  x"cb",  x"10",  x"cb",  x"21",  x"cb",  x"10", -- 0838
         x"ed",  x"b8",  x"23",  x"18",  x"b1",  x"2a",  x"1a",  x"00", -- 0840
         x"ed",  x"4b",  x"1e",  x"00",  x"b7",  x"ed",  x"42",  x"c8", -- 0848
         x"cd",  x"05",  x"d7",  x"d8",  x"11",  x"16",  x"00",  x"cd", -- 0850
         x"4a",  x"d6",  x"2a",  x"1a",  x"00",  x"ed",  x"5b",  x"1e", -- 0858
         x"00",  x"ed",  x"52",  x"cc",  x"be",  x"d2",  x"18",  x"15", -- 0860
         x"2a",  x"1c",  x"00",  x"ed",  x"4b",  x"18",  x"00",  x"b7", -- 0868
         x"ed",  x"42",  x"c8",  x"cd",  x"05",  x"d7",  x"d8",  x"11", -- 0870
         x"16",  x"00",  x"cd",  x"9f",  x"d6",  x"cd",  x"f0",  x"d7", -- 0878
         x"c3",  x"e4",  x"c6",  x"2a",  x"9c",  x"b7",  x"cd",  x"89", -- 0880
         x"c5",  x"54",  x"5d",  x"13",  x"3a",  x"9f",  x"b7",  x"87", -- 0888
         x"4f",  x"87",  x"87",  x"81",  x"3d",  x"06",  x"00",  x"4f", -- 0890
         x"3a",  x"9e",  x"b7",  x"cb",  x"3f",  x"e5",  x"d5",  x"c5", -- 0898
         x"36",  x"00",  x"ed",  x"b0",  x"c1",  x"d1",  x"e1",  x"24", -- 08A0
         x"14",  x"3d",  x"20",  x"f1",  x"ed",  x"4b",  x"9e",  x"b7", -- 08A8
         x"50",  x"cd",  x"03",  x"f0",  x"41",  x"4f",  x"ed",  x"5b", -- 08B0
         x"9c",  x"b7",  x"cd",  x"60",  x"c5",  x"54",  x"5d",  x"13", -- 08B8
         x"0b",  x"36",  x"00",  x"ed",  x"b0",  x"16",  x"00",  x"1e", -- 08C0
         x"00",  x"c9",  x"ed",  x"5b",  x"9e",  x"b7",  x"15",  x"1d", -- 08C8
         x"c9",  x"7b",  x"a7",  x"28",  x"03",  x"1d",  x"18",  x"0f", -- 08D0
         x"7a",  x"a7",  x"20",  x"05",  x"cd",  x"42",  x"c7",  x"d8", -- 08D8
         x"3e",  x"15",  x"3a",  x"9e",  x"b7",  x"3d",  x"5f",  x"7b", -- 08E0
         x"e6",  x"07",  x"c8",  x"cd",  x"60",  x"c5",  x"7e",  x"b7", -- 08E8
         x"c0",  x"2b",  x"7e",  x"b7",  x"28",  x"db",  x"c9",  x"cd", -- 08F0
         x"d1",  x"c8",  x"d8",  x"cd",  x"60",  x"c5",  x"7e",  x"fe", -- 08F8
         x"21",  x"30",  x"f4",  x"cd",  x"60",  x"c5",  x"7e",  x"fe", -- 0900
         x"21",  x"30",  x"0d",  x"cd",  x"d1",  x"c8",  x"d8",  x"18", -- 0908
         x"f2",  x"cd",  x"d1",  x"c8",  x"d8",  x"cd",  x"60",  x"c5", -- 0910
         x"2b",  x"7e",  x"fe",  x"21",  x"d8",  x"18",  x"f2",  x"d5", -- 0918
         x"cd",  x"96",  x"ca",  x"2a",  x"99",  x"b7",  x"cd",  x"30", -- 0920
         x"c9",  x"cd",  x"37",  x"ca",  x"d1",  x"c3",  x"6e",  x"d9", -- 0928
         x"e9",  x"21",  x"3e",  x"00",  x"7e",  x"c6",  x"20",  x"77", -- 0930
         x"e6",  x"60",  x"fe",  x"60",  x"28",  x"f6",  x"11",  x"00", -- 0938
         x"00",  x"21",  x"a0",  x"ad",  x"7e",  x"23",  x"fe",  x"40", -- 0940
         x"28",  x"14",  x"fe",  x"60",  x"28",  x"10",  x"fe",  x"5b", -- 0948
         x"38",  x"0f",  x"fe",  x"5e",  x"38",  x"08",  x"fe",  x"7b", -- 0950
         x"38",  x"07",  x"fe",  x"7f",  x"30",  x"03",  x"cd",  x"b4", -- 0958
         x"c5",  x"1c",  x"3e",  x"50",  x"93",  x"20",  x"dd",  x"5f", -- 0960
         x"14",  x"3e",  x"17",  x"ba",  x"20",  x"d6",  x"18",  x"12", -- 0968
         x"3a",  x"3e",  x"00",  x"ee",  x"10",  x"32",  x"3e",  x"00", -- 0970
         x"18",  x"08",  x"dd",  x"7e",  x"08",  x"ee",  x"20",  x"dd", -- 0978
         x"77",  x"08",  x"cd",  x"40",  x"d8",  x"ed",  x"5b",  x"20", -- 0980
         x"00",  x"ed",  x"53",  x"a0",  x"b7",  x"c9",  x"7b",  x"a7", -- 0988
         x"28",  x"03",  x"1d",  x"18",  x"10",  x"7a",  x"a7",  x"20", -- 0990
         x"09",  x"3c",  x"32",  x"a1",  x"b7",  x"cd",  x"42",  x"c7", -- 0998
         x"d8",  x"3e",  x"15",  x"1e",  x"4f",  x"cd",  x"60",  x"c5", -- 09A0
         x"7e",  x"a7",  x"20",  x"10",  x"7d",  x"e6",  x"f8",  x"6f", -- 09A8
         x"7e",  x"a7",  x"20",  x"02",  x"36",  x"20",  x"23",  x"7d", -- 09B0
         x"e6",  x"07",  x"20",  x"f4",  x"ed",  x"5b",  x"a0",  x"b7", -- 09B8
         x"cd",  x"d1",  x"c8",  x"d8",  x"d5",  x"cd",  x"60",  x"c5", -- 09C0
         x"7e",  x"b7",  x"28",  x"24",  x"e5",  x"d5",  x"1c",  x"cd", -- 09C8
         x"60",  x"c5",  x"30",  x"08",  x"1e",  x"00",  x"14",  x"cd", -- 09D0
         x"60",  x"c5",  x"38",  x"0f",  x"7e",  x"a7",  x"28",  x"0b", -- 09D8
         x"42",  x"4b",  x"d1",  x"e3",  x"cd",  x"b1",  x"c5",  x"50", -- 09E0
         x"59",  x"18",  x"e2",  x"d1",  x"e1",  x"cd",  x"b0",  x"c5", -- 09E8
         x"d1",  x"c9",  x"f5",  x"db",  x"88",  x"e6",  x"5b",  x"d3", -- 09F0
         x"88",  x"f1",  x"c9",  x"cd",  x"5a",  x"00",  x"ed",  x"b0", -- 09F8
         x"18",  x"2c",  x"cd",  x"5a",  x"00",  x"ed",  x"b8",  x"18", -- 0A00
         x"25",  x"cd",  x"5a",  x"00",  x"ed",  x"b1",  x"18",  x"1e", -- 0A08
         x"cd",  x"5a",  x"00",  x"ed",  x"b9",  x"18",  x"17",  x"cd", -- 0A10
         x"5a",  x"00",  x"ed",  x"a1",  x"18",  x"10",  x"cd",  x"5a", -- 0A18
         x"00",  x"7e",  x"18",  x"0a",  x"cd",  x"5a",  x"00",  x"0a", -- 0A20
         x"18",  x"04",  x"cd",  x"5a",  x"00",  x"77",  x"f5",  x"db", -- 0A28
         x"88",  x"f6",  x"a4",  x"d3",  x"88",  x"f1",  x"c9",  x"2a", -- 0A30
         x"b0",  x"b7",  x"5e",  x"23",  x"56",  x"ed",  x"53",  x"d0", -- 0A38
         x"b4",  x"11",  x"36",  x"c6",  x"72",  x"2b",  x"73",  x"11", -- 0A40
         x"4a",  x"00",  x"19",  x"5e",  x"23",  x"56",  x"ed",  x"53", -- 0A48
         x"d2",  x"b4",  x"11",  x"43",  x"c6",  x"72",  x"2b",  x"73", -- 0A50
         x"2a",  x"dd",  x"b7",  x"22",  x"d4",  x"b4",  x"3a",  x"df", -- 0A58
         x"b7",  x"32",  x"d6",  x"b4",  x"21",  x"eb",  x"b4",  x"22", -- 0A60
         x"dd",  x"b7",  x"3e",  x"24",  x"32",  x"df",  x"b7",  x"11", -- 0A68
         x"5d",  x"db",  x"06",  x"0a",  x"73",  x"23",  x"72",  x"23", -- 0A70
         x"10",  x"fa",  x"eb",  x"21",  x"54",  x"df",  x"01",  x"34", -- 0A78
         x"00",  x"ed",  x"b0",  x"21",  x"20",  x"00",  x"22",  x"de", -- 0A80
         x"b4",  x"21",  x"00",  x"00",  x"22",  x"9c",  x"b7",  x"21", -- 0A88
         x"50",  x"19",  x"22",  x"9e",  x"b7",  x"c9",  x"2a",  x"b0", -- 0A90
         x"b7",  x"ed",  x"5b",  x"d0",  x"b4",  x"73",  x"23",  x"72", -- 0A98
         x"11",  x"49",  x"00",  x"19",  x"ed",  x"5b",  x"d2",  x"b4", -- 0AA0
         x"73",  x"23",  x"72",  x"2a",  x"d4",  x"b4",  x"22",  x"dd", -- 0AA8
         x"b7",  x"3a",  x"d6",  x"b4",  x"32",  x"df",  x"b7",  x"21", -- 0AB0
         x"00",  x"00",  x"22",  x"9c",  x"b7",  x"21",  x"28",  x"20", -- 0AB8
         x"22",  x"9e",  x"b7",  x"cd",  x"03",  x"f0",  x"20",  x"3e", -- 0AC0
         x"12",  x"cd",  x"03",  x"f0",  x"00",  x"c9",  x"06",  x"08", -- 0AC8
         x"0e",  x"80",  x"ed",  x"78",  x"fe",  x"f6",  x"28",  x"09", -- 0AD0
         x"fe",  x"f4",  x"28",  x"05",  x"04",  x"20",  x"f1",  x"18", -- 0AD8
         x"09",  x"16",  x"c3",  x"68",  x"3e",  x"02",  x"cd",  x"03", -- 0AE0
         x"f0",  x"26",  x"21",  x"f2",  x"c9",  x"11",  x"5a",  x"00", -- 0AE8
         x"01",  x"45",  x"00",  x"ed",  x"b0",  x"c9",  x"7f",  x"7f", -- 0AF0
         x"45",  x"44",  x"49",  x"54",  x"01",  x"32",  x"e7",  x"bf", -- 0AF8
         x"cd",  x"e5",  x"d1",  x"cd",  x"ce",  x"ca",  x"21",  x"00", -- 0B00
         x"02",  x"36",  x"0d",  x"23",  x"22",  x"18",  x"00",  x"22", -- 0B08
         x"1c",  x"00",  x"23",  x"2e",  x"ff",  x"cd",  x"86",  x"00", -- 0B10
         x"4f",  x"2f",  x"cd",  x"92",  x"00",  x"cd",  x"86",  x"00", -- 0B18
         x"2f",  x"b9",  x"79",  x"cd",  x"92",  x"00",  x"20",  x"03", -- 0B20
         x"24",  x"18",  x"ea",  x"25",  x"3e",  x"03",  x"cd",  x"92", -- 0B28
         x"00",  x"22",  x"1a",  x"00",  x"22",  x"1e",  x"00",  x"21", -- 0B30
         x"00",  x"00",  x"22",  x"20",  x"00",  x"cd",  x"d7",  x"cd", -- 0B38
         x"af",  x"32",  x"22",  x"00",  x"21",  x"08",  x"48",  x"22", -- 0B40
         x"10",  x"00",  x"18",  x"0c",  x"7f",  x"7f",  x"52",  x"45", -- 0B48
         x"45",  x"44",  x"49",  x"54",  x"01",  x"cd",  x"ce",  x"ca", -- 0B50
         x"01",  x"f1",  x"83",  x"ed",  x"79",  x"cd",  x"b7",  x"ca", -- 0B58
         x"cd",  x"03",  x"f0",  x"23",  x"0c",  x"00",  x"21",  x"a2", -- 0B60
         x"b7",  x"cb",  x"ce",  x"21",  x"3e",  x"00",  x"36",  x"00", -- 0B68
         x"01",  x"80",  x"fc",  x"ed",  x"78",  x"fe",  x"a7",  x"20", -- 0B70
         x"0d",  x"34",  x"01",  x"f1",  x"83",  x"ed",  x"78",  x"3c", -- 0B78
         x"fe",  x"21",  x"38",  x"02",  x"cb",  x"ce",  x"21",  x"00", -- 0B80
         x"00",  x"06",  x"ff",  x"7e",  x"23",  x"fe",  x"7f",  x"28", -- 0B88
         x"04",  x"fe",  x"dd",  x"20",  x"05",  x"be",  x"20",  x"02", -- 0B90
         x"36",  x"00",  x"10",  x"ef",  x"01",  x"d1",  x"18",  x"18", -- 0B98
         x"0b",  x"dd",  x"dd",  x"4d",  x"45",  x"4e",  x"55",  x"1f", -- 0BA0
         x"e1",  x"01",  x"00",  x"47",  x"c5",  x"cd",  x"b7",  x"ca", -- 0BA8
         x"cd",  x"03",  x"f0",  x"23",  x"0c",  x"0a",  x"0a",  x"00", -- 0BB0
         x"06",  x"28",  x"cd",  x"03",  x"f0",  x"23",  x"5f",  x"00", -- 0BB8
         x"10",  x"f8",  x"cd",  x"63",  x"cc",  x"cd",  x"e7",  x"cc", -- 0BC0
         x"cd",  x"ae",  x"cc",  x"cd",  x"03",  x"f0",  x"2d",  x"21", -- 0BC8
         x"00",  x"ba",  x"c1",  x"cd",  x"03",  x"f0",  x"23",  x"02", -- 0BD0
         x"2d",  x"00",  x"cd",  x"03",  x"f0",  x"2a",  x"38",  x"4a", -- 0BD8
         x"3e",  x"dd",  x"ed",  x"b1",  x"e2",  x"2a",  x"cc",  x"ed", -- 0BE0
         x"a1",  x"20",  x"f7",  x"7e",  x"fe",  x"20",  x"38",  x"0f", -- 0BE8
         x"fe",  x"30",  x"38",  x"df",  x"fe",  x"5f",  x"30",  x"db", -- 0BF0
         x"cd",  x"8c",  x"ce",  x"23",  x"0b",  x"18",  x"ec",  x"cd", -- 0BF8
         x"87",  x"ce",  x"18",  x"cf",  x"e1",  x"cd",  x"ea",  x"de", -- 0C00
         x"18",  x"06",  x"3e",  x"0b",  x"cd",  x"03",  x"f0",  x"00", -- 0C08
         x"3e",  x"02",  x"cd",  x"03",  x"f0",  x"00",  x"cd",  x"03", -- 0C10
         x"f0",  x"20",  x"cd",  x"63",  x"cc",  x"cd",  x"ae",  x"cc", -- 0C18
         x"cd",  x"e7",  x"cc",  x"cd",  x"03",  x"f0",  x"23",  x"0d", -- 0C20
         x"2d",  x"00",  x"cd",  x"03",  x"f0",  x"17",  x"38",  x"da", -- 0C28
         x"13",  x"1a",  x"fe",  x"20",  x"28",  x"ed",  x"a7",  x"28", -- 0C30
         x"ea",  x"3e",  x"dd",  x"21",  x"00",  x"ba",  x"01",  x"00", -- 0C38
         x"47",  x"cd",  x"03",  x"f0",  x"1d",  x"30",  x"be",  x"7e", -- 0C40
         x"23",  x"e5",  x"fe",  x"1f",  x"28",  x"10",  x"cd",  x"03", -- 0C48
         x"f0",  x"22",  x"38",  x"b0",  x"21",  x"16",  x"cc",  x"e3", -- 0C50
         x"e5",  x"cd",  x"03",  x"f0",  x"15",  x"c9",  x"21",  x"16", -- 0C58
         x"cc",  x"e3",  x"e9",  x"2a",  x"a0",  x"b7",  x"e5",  x"cd", -- 0C60
         x"b7",  x"ca",  x"21",  x"01",  x"01",  x"22",  x"a0",  x"b7", -- 0C68
         x"21",  x"f5",  x"b7",  x"7e",  x"fe",  x"21",  x"38",  x"1c", -- 0C70
         x"cd",  x"03",  x"f0",  x"23",  x"45",  x"44",  x"49",  x"54", -- 0C78
         x"3a",  x"00",  x"06",  x"08",  x"cd",  x"2b",  x"d6",  x"3e", -- 0C80
         x"2e",  x"cd",  x"03",  x"f0",  x"00",  x"06",  x"03",  x"cd", -- 0C88
         x"2b",  x"d6",  x"18",  x"42",  x"cd",  x"03",  x"f0",  x"23", -- 0C90
         x"3e",  x"3e",  x"20",  x"4b",  x"43",  x"2d",  x"45",  x"44", -- 0C98
         x"49",  x"54",  x"20",  x"30",  x"2e",  x"34",  x"20",  x"3c", -- 0CA0
         x"3c",  x"0d",  x"0a",  x"00",  x"18",  x"28",  x"2a",  x"a0", -- 0CA8
         x"b7",  x"e5",  x"cd",  x"b7",  x"ca",  x"21",  x"1d",  x"01", -- 0CB0
         x"22",  x"a0",  x"b7",  x"cd",  x"03",  x"f0",  x"23",  x"46", -- 0CB8
         x"72",  x"65",  x"69",  x"3a",  x"1f",  x"1f",  x"1f",  x"1f", -- 0CC0
         x"00",  x"2a",  x"1e",  x"00",  x"ed",  x"5b",  x"1c",  x"00", -- 0CC8
         x"af",  x"ed",  x"52",  x"cd",  x"f6",  x"de",  x"e1",  x"22", -- 0CD0
         x"a0",  x"b7",  x"21",  x"00",  x"04",  x"22",  x"9c",  x"b7", -- 0CD8
         x"21",  x"28",  x"1c",  x"22",  x"9e",  x"b7",  x"c9",  x"2a", -- 0CE0
         x"a0",  x"b7",  x"e5",  x"cd",  x"b7",  x"ca",  x"21",  x"13", -- 0CE8
         x"01",  x"22",  x"a0",  x"b7",  x"3e",  x"28",  x"cd",  x"03", -- 0CF0
         x"f0",  x"00",  x"06",  x"09",  x"cd",  x"03",  x"f0",  x"2b", -- 0CF8
         x"10",  x"fa",  x"3e",  x"14",  x"32",  x"a0",  x"b7",  x"3e", -- 0D00
         x"fe",  x"cd",  x"03",  x"f0",  x"49",  x"11",  x"14",  x"01", -- 0D08
         x"cd",  x"03",  x"f0",  x"32",  x"11",  x"53",  x"cd",  x"01", -- 0D10
         x"04",  x"00",  x"1a",  x"13",  x"ed",  x"a1",  x"20",  x"2b", -- 0D18
         x"ea",  x"1a",  x"cd",  x"21",  x"3e",  x"00",  x"cb",  x"4e", -- 0D20
         x"28",  x"21",  x"cd",  x"03",  x"f0",  x"23",  x"3a",  x"00", -- 0D28
         x"3e",  x"01",  x"01",  x"f1",  x"80",  x"ed",  x"79",  x"ed", -- 0D30
         x"78",  x"cb",  x"47",  x"20",  x"fa",  x"04",  x"ed",  x"78", -- 0D38
         x"cd",  x"8c",  x"ce",  x"04",  x"ed",  x"68",  x"26",  x"00", -- 0D40
         x"cd",  x"f6",  x"de",  x"3e",  x"29",  x"cd",  x"03",  x"f0", -- 0D48
         x"00",  x"18",  x"83",  x"44",  x"49",  x"53",  x"4b",  x"dd", -- 0D50
         x"dd",  x"51",  x"55",  x"49",  x"54",  x"1f",  x"cd",  x"b7", -- 0D58
         x"ca",  x"21",  x"a1",  x"b7",  x"7e",  x"c6",  x"04",  x"77", -- 0D60
         x"23",  x"cb",  x"8e",  x"11",  x"89",  x"cd",  x"21",  x"00", -- 0D68
         x"e0",  x"01",  x"00",  x"20",  x"dd",  x"7e",  x"09",  x"cd", -- 0D70
         x"03",  x"f0",  x"1d",  x"23",  x"e3",  x"ed",  x"5b",  x"7f", -- 0D78
         x"b7",  x"3e",  x"02",  x"6f",  x"1e",  x"26",  x"c3",  x"09", -- 0D80
         x"f0",  x"4d",  x"45",  x"4e",  x"55",  x"00",  x"dd",  x"dd", -- 0D88
         x"43",  x"4c",  x"45",  x"41",  x"52",  x"1f",  x"2a",  x"1c", -- 0D90
         x"00",  x"ed",  x"5b",  x"18",  x"00",  x"a7",  x"ed",  x"52", -- 0D98
         x"44",  x"4d",  x"2a",  x"1a",  x"00",  x"ed",  x"5b",  x"1e", -- 0DA0
         x"00",  x"ed",  x"52",  x"09",  x"7c",  x"b5",  x"28",  x"27", -- 0DA8
         x"cd",  x"03",  x"f0",  x"23",  x"0d",  x"44",  x"65",  x"6c", -- 0DB0
         x"65",  x"74",  x"65",  x"20",  x"54",  x"65",  x"78",  x"74", -- 0DB8
         x"00",  x"cd",  x"65",  x"d5",  x"d8",  x"2a",  x"18",  x"00", -- 0DC0
         x"22",  x"1c",  x"00",  x"2a",  x"1a",  x"00",  x"22",  x"1e", -- 0DC8
         x"00",  x"cd",  x"ae",  x"cc",  x"cd",  x"e2",  x"cd",  x"21", -- 0DD0
         x"f5",  x"b7",  x"06",  x"0b",  x"36",  x"20",  x"23",  x"10", -- 0DD8
         x"fb",  x"c9",  x"11",  x"00",  x"00",  x"ed",  x"53",  x"20", -- 0DE0
         x"00",  x"c9",  x"dd",  x"dd",  x"53",  x"41",  x"56",  x"45", -- 0DE8
         x"1f",  x"cd",  x"9c",  x"d6",  x"ed",  x"5b",  x"1e",  x"00", -- 0DF0
         x"2a",  x"1a",  x"00",  x"af",  x"ed",  x"52",  x"c8",  x"cd", -- 0DF8
         x"f0",  x"d5",  x"d8",  x"cd",  x"87",  x"ce",  x"cd",  x"36", -- 0E00
         x"d6",  x"ed",  x"5b",  x"1e",  x"00",  x"dd",  x"36",  x"02", -- 0E08
         x"01",  x"dd",  x"cb",  x"07",  x"fe",  x"3e",  x"08",  x"cd", -- 0E10
         x"03",  x"f0",  x"49",  x"28",  x"18",  x"21",  x"80",  x"b7", -- 0E18
         x"45",  x"3e",  x"1a",  x"2d",  x"77",  x"20",  x"fc",  x"eb", -- 0E20
         x"cd",  x"86",  x"00",  x"eb",  x"13",  x"77",  x"fe",  x"03", -- 0E28
         x"28",  x"03",  x"23",  x"10",  x"f2",  x"dd",  x"7e",  x"02", -- 0E30
         x"cd",  x"03",  x"f0",  x"1c",  x"cd",  x"03",  x"f0",  x"23", -- 0E38
         x"08",  x"08",  x"00",  x"cd",  x"03",  x"f0",  x"2a",  x"01", -- 0E40
         x"a0",  x"00",  x"38",  x"23",  x"2a",  x"1a",  x"00",  x"ed", -- 0E48
         x"52",  x"38",  x"1c",  x"d5",  x"dd",  x"cb",  x"07",  x"7e", -- 0E50
         x"28",  x"0d",  x"dd",  x"cb",  x"07",  x"be",  x"21",  x"00", -- 0E58
         x"00",  x"cd",  x"03",  x"f0",  x"08",  x"18",  x"04",  x"cd", -- 0E60
         x"03",  x"f0",  x"01",  x"d1",  x"d8",  x"18",  x"ae",  x"dd", -- 0E68
         x"cb",  x"07",  x"7e",  x"28",  x"0b",  x"dd",  x"cb",  x"07", -- 0E70
         x"be",  x"21",  x"00",  x"00",  x"cd",  x"03",  x"f0",  x"08", -- 0E78
         x"cd",  x"03",  x"f0",  x"09",  x"d4",  x"59",  x"cf",  x"cd", -- 0E80
         x"03",  x"f0",  x"2c",  x"c9",  x"cd",  x"03",  x"f0",  x"24", -- 0E88
         x"c9",  x"dd",  x"dd",  x"4c",  x"4f",  x"41",  x"44",  x"1f", -- 0E90
         x"3e",  x"08",  x"cd",  x"03",  x"f0",  x"49",  x"28",  x"07", -- 0E98
         x"cd",  x"f0",  x"d5",  x"d8",  x"cd",  x"87",  x"ce",  x"cd", -- 0EA0
         x"e2",  x"cd",  x"21",  x"00",  x"b7",  x"dd",  x"75",  x"05", -- 0EA8
         x"dd",  x"74",  x"06",  x"dd",  x"cb",  x"07",  x"c6",  x"21", -- 0EB0
         x"00",  x"00",  x"cd",  x"03",  x"f0",  x"0a",  x"d8",  x"af", -- 0EB8
         x"cd",  x"65",  x"cf",  x"da",  x"29",  x"cf",  x"3e",  x"08", -- 0EC0
         x"cd",  x"03",  x"f0",  x"49",  x"20",  x"1c",  x"3e",  x"02", -- 0EC8
         x"cd",  x"8c",  x"ce",  x"11",  x"00",  x"00",  x"21",  x"00", -- 0ED0
         x"b7",  x"01",  x"0b",  x"00",  x"7e",  x"fe",  x"20",  x"d4", -- 0ED8
         x"8c",  x"ce",  x"ed",  x"a0",  x"ea",  x"dc",  x"ce",  x"cd", -- 0EE0
         x"87",  x"ce",  x"dd",  x"36",  x"03",  x"02",  x"ed",  x"5b", -- 0EE8
         x"1c",  x"00",  x"2a",  x"1e",  x"00",  x"af",  x"ed",  x"52", -- 0EF0
         x"28",  x"2b",  x"e5",  x"cd",  x"65",  x"cf",  x"e1",  x"38", -- 0EF8
         x"28",  x"01",  x"80",  x"00",  x"ed",  x"42",  x"30",  x"02", -- 0F00
         x"09",  x"4d",  x"41",  x"21",  x"00",  x"b7",  x"7e",  x"fe", -- 0F08
         x"03",  x"28",  x"16",  x"fe",  x"1a",  x"28",  x"12",  x"23", -- 0F10
         x"eb",  x"cd",  x"92",  x"00",  x"eb",  x"13",  x"10",  x"ee", -- 0F18
         x"dd",  x"34",  x"03",  x"18",  x"cd",  x"3c",  x"32",  x"22", -- 0F20
         x"00",  x"cd",  x"03",  x"f0",  x"0b",  x"62",  x"6b",  x"ed", -- 0F28
         x"4b",  x"1c",  x"00",  x"a7",  x"ed",  x"42",  x"ca",  x"87", -- 0F30
         x"ce",  x"44",  x"4d",  x"2a",  x"1e",  x"00",  x"eb",  x"cd", -- 0F38
         x"87",  x"ce",  x"1b",  x"2b",  x"cd",  x"6a",  x"00",  x"13", -- 0F40
         x"23",  x"ed",  x"53",  x"1e",  x"00",  x"3a",  x"22",  x"00", -- 0F48
         x"b7",  x"28",  x"06",  x"cd",  x"41",  x"d5",  x"c3",  x"87", -- 0F50
         x"ce",  x"21",  x"00",  x"00",  x"11",  x"f5",  x"b7",  x"01", -- 0F58
         x"0b",  x"00",  x"ed",  x"b0",  x"c9",  x"2e",  x"04",  x"20", -- 0F60
         x"06",  x"dd",  x"cb",  x"07",  x"fe",  x"18",  x"35",  x"cd", -- 0F68
         x"03",  x"f0",  x"2a",  x"d8",  x"dd",  x"7e",  x"03",  x"fe", -- 0F70
         x"02",  x"20",  x"24",  x"dd",  x"cb",  x"07",  x"7e",  x"28", -- 0F78
         x"1e",  x"dd",  x"cb",  x"07",  x"be",  x"d9",  x"ed",  x"4b", -- 0F80
         x"11",  x"b7",  x"2a",  x"13",  x"b7",  x"ed",  x"42",  x"22", -- 0F88
         x"86",  x"b7",  x"d9",  x"3a",  x"10",  x"b7",  x"fe",  x"03", -- 0F90
         x"38",  x"05",  x"dd",  x"35",  x"03",  x"18",  x"05",  x"cd", -- 0F98
         x"03",  x"f0",  x"05",  x"d8",  x"3e",  x"01",  x"3d",  x"dd", -- 0FA0
         x"7e",  x"02",  x"f5",  x"dd",  x"be",  x"03",  x"28",  x"08", -- 0FA8
         x"3c",  x"20",  x"21",  x"7d",  x"fe",  x"04",  x"20",  x"1c", -- 0FB0
         x"f1",  x"38",  x"08",  x"f5",  x"3e",  x"02",  x"cd",  x"03", -- 0FB8
         x"f0",  x"00",  x"f1",  x"f5",  x"cd",  x"03",  x"f0",  x"1c", -- 0FC0
         x"f1",  x"38",  x"0f",  x"cd",  x"03",  x"f0",  x"23",  x"3e", -- 0FC8
         x"20",  x"00",  x"a7",  x"c9",  x"f1",  x"37",  x"2c",  x"2d", -- 0FD0
         x"18",  x"e9",  x"28",  x"0b",  x"cd",  x"03",  x"f0",  x"23", -- 0FD8
         x"2a",  x"08",  x"08",  x"08",  x"00",  x"18",  x"88",  x"67", -- 0FE0
         x"2d",  x"28",  x"0b",  x"cd",  x"03",  x"f0",  x"23",  x"3f", -- 0FE8
         x"20",  x"07",  x"00",  x"c3",  x"6f",  x"cf",  x"cd",  x"03", -- 0FF0
         x"f0",  x"23",  x"21",  x"0a",  x"0d",  x"00",  x"a7",  x"c9", -- 0FF8
         x"dd",  x"dd",  x"50",  x"52",  x"49",  x"4e",  x"54",  x"01", -- 1000
         x"cd",  x"e9",  x"d0",  x"d8",  x"cd",  x"9c",  x"d6",  x"2a", -- 1008
         x"1e",  x"00",  x"1e",  x"00",  x"3a",  x"82",  x"b7",  x"47", -- 1010
         x"cd",  x"86",  x"00",  x"23",  x"fe",  x"03",  x"28",  x"7d", -- 1018
         x"fe",  x"0d",  x"20",  x"11",  x"cd",  x"ab",  x"d0",  x"38", -- 1020
         x"7d",  x"04",  x"05",  x"28",  x"eb",  x"10",  x"e9",  x"3a", -- 1028
         x"82",  x"b7",  x"47",  x"3e",  x"0c",  x"fe",  x"0e",  x"28", -- 1030
         x"4e",  x"fe",  x"0f",  x"20",  x"42",  x"cd",  x"86",  x"00", -- 1038
         x"fe",  x"20",  x"20",  x"03",  x"23",  x"18",  x"f6",  x"d5", -- 1040
         x"e5",  x"11",  x"80",  x"a8",  x"cd",  x"86",  x"00",  x"fe", -- 1048
         x"21",  x"38",  x"05",  x"12",  x"13",  x"23",  x"18",  x"f4", -- 1050
         x"af",  x"12",  x"11",  x"80",  x"a8",  x"e5",  x"cd",  x"03", -- 1058
         x"f0",  x"18",  x"e1",  x"30",  x"04",  x"e1",  x"d1",  x"18", -- 1060
         x"1e",  x"d1",  x"d1",  x"3a",  x"97",  x"b7",  x"cd",  x"8c", -- 1068
         x"ce",  x"cd",  x"86",  x"00",  x"23",  x"fe",  x"0d",  x"28", -- 1070
         x"1c",  x"fe",  x"03",  x"28",  x"20",  x"18",  x"c8",  x"1c", -- 1078
         x"1d",  x"20",  x"12",  x"fe",  x"2e",  x"20",  x"0e",  x"cd", -- 1080
         x"86",  x"00",  x"23",  x"fe",  x"03",  x"28",  x"0e",  x"fe", -- 1088
         x"0a",  x"20",  x"f4",  x"18",  x"83",  x"cd",  x"ab",  x"d0", -- 1090
         x"38",  x"0c",  x"c3",  x"18",  x"d0",  x"3a",  x"82",  x"b7", -- 1098
         x"b8",  x"3e",  x"0c",  x"c4",  x"ab",  x"d0",  x"cd",  x"03", -- 10A0
         x"f0",  x"20",  x"c9",  x"c5",  x"06",  x"01",  x"fe",  x"20", -- 10A8
         x"30",  x"21",  x"fe",  x"0c",  x"28",  x"09",  x"fe",  x"0d", -- 10B0
         x"20",  x"09",  x"cd",  x"8c",  x"ce",  x"3e",  x"0a",  x"1e", -- 10B8
         x"ff",  x"18",  x"10",  x"fe",  x"09",  x"20",  x"14",  x"3e", -- 10C0
         x"08",  x"93",  x"e6",  x"07",  x"20",  x"02",  x"3e",  x"08", -- 10C8
         x"47",  x"3e",  x"20",  x"cd",  x"8c",  x"ce",  x"1c",  x"10", -- 10D0
         x"fa",  x"18",  x"09",  x"d6",  x"10",  x"38",  x"05",  x"fe", -- 10D8
         x"0a",  x"dc",  x"60",  x"d1",  x"cd",  x"da",  x"d4",  x"c1", -- 10E0
         x"c9",  x"2a",  x"be",  x"b7",  x"7e",  x"fe",  x"c9",  x"20", -- 10E8
         x"1c",  x"cd",  x"03",  x"f0",  x"23",  x"4b",  x"65",  x"69", -- 10F0
         x"6e",  x"20",  x"44",  x"72",  x"75",  x"63",  x"6b",  x"65", -- 10F8
         x"72",  x"20",  x"61",  x"6b",  x"74",  x"69",  x"76",  x"21", -- 1100
         x"0d",  x"0a",  x"00",  x"37",  x"c9",  x"3a",  x"81",  x"b7", -- 1108
         x"b7",  x"28",  x"20",  x"3a",  x"82",  x"b7",  x"e6",  x"f0", -- 1110
         x"0f",  x"0f",  x"0f",  x"0f",  x"fe",  x"0a",  x"30",  x"28", -- 1118
         x"3c",  x"47",  x"3e",  x"f6",  x"c6",  x"0a",  x"10",  x"fc", -- 1120
         x"47",  x"3a",  x"82",  x"b7",  x"e6",  x"0f",  x"fe",  x"0a", -- 1128
         x"30",  x"16",  x"80",  x"32",  x"82",  x"b7",  x"21",  x"08", -- 1130
         x"f0",  x"cd",  x"03",  x"f0",  x"1e",  x"21",  x"e1",  x"b4", -- 1138
         x"af",  x"06",  x"0a",  x"77",  x"23",  x"10",  x"fc",  x"c9", -- 1140
         x"cd",  x"03",  x"f0",  x"23",  x"50",  x"61",  x"72",  x"61", -- 1148
         x"6d",  x"65",  x"74",  x"65",  x"72",  x"66",  x"65",  x"68", -- 1150
         x"6c",  x"65",  x"72",  x"0d",  x"0a",  x"00",  x"37",  x"c9", -- 1158
         x"e5",  x"21",  x"e1",  x"b4",  x"06",  x"00",  x"4f",  x"09", -- 1160
         x"7e",  x"ee",  x"01",  x"77",  x"81",  x"81",  x"4f",  x"0c", -- 1168
         x"21",  x"86",  x"d1",  x"46",  x"23",  x"0d",  x"28",  x"05", -- 1170
         x"23",  x"10",  x"fd",  x"18",  x"f6",  x"7e",  x"cd",  x"8c", -- 1178
         x"ce",  x"23",  x"10",  x"f9",  x"e1",  x"c9",  x"03",  x"1b", -- 1180
         x"55",  x"00",  x"03",  x"1b",  x"55",  x"01",  x"02",  x"1b", -- 1188
         x"54",  x"03",  x"1b",  x"53",  x"00",  x"01",  x"12",  x"01", -- 1190
         x"0f",  x"03",  x"1b",  x"2d",  x"30",  x"03",  x"1b",  x"2d", -- 1198
         x"31",  x"02",  x"1b",  x"50",  x"02",  x"1b",  x"4d",  x"03", -- 11A0
         x"1b",  x"57",  x"00",  x"03",  x"1b",  x"57",  x"01",  x"02", -- 11A8
         x"1b",  x"48",  x"02",  x"1b",  x"47",  x"02",  x"1b",  x"54", -- 11B0
         x"03",  x"1b",  x"53",  x"01",  x"02",  x"1b",  x"46",  x"02", -- 11B8
         x"1b",  x"45",  x"03",  x"1b",  x"78",  x"00",  x"03",  x"1b", -- 11C0
         x"78",  x"01",  x"dd",  x"dd",  x"4b",  x"45",  x"59",  x"01", -- 11C8
         x"b7",  x"20",  x"05",  x"cd",  x"03",  x"f0",  x"3a",  x"c9", -- 11D0
         x"7d",  x"b7",  x"28",  x"09",  x"fe",  x"d5",  x"28",  x"0c", -- 11D8
         x"cd",  x"03",  x"f0",  x"39",  x"c9",  x"21",  x"11",  x"d2", -- 11E0
         x"06",  x"03",  x"18",  x"05",  x"21",  x"06",  x"d2",  x"06", -- 11E8
         x"0b",  x"11",  x"00",  x"b9",  x"af",  x"12",  x"13",  x"ed", -- 11F0
         x"a0",  x"03",  x"10",  x"f9",  x"eb",  x"36",  x"00",  x"23", -- 11F8
         x"7d",  x"fe",  x"9c",  x"20",  x"f8",  x"c9",  x"5b",  x"5c", -- 1200
         x"5d",  x"7e",  x"05",  x"06",  x"7b",  x"7c",  x"7d",  x"60", -- 1208
         x"7f",  x"1b",  x"05",  x"06",  x"3a",  x"21",  x"00",  x"16", -- 1210
         x"00",  x"5f",  x"b7",  x"c4",  x"4a",  x"d6",  x"cd",  x"e2", -- 1218
         x"cd",  x"ed",  x"5b",  x"1e",  x"00",  x"2a",  x"1a",  x"00", -- 1220
         x"af",  x"ed",  x"52",  x"ca",  x"b8",  x"d2",  x"44",  x"4d", -- 1228
         x"eb",  x"11",  x"23",  x"00",  x"1a",  x"b7",  x"c8",  x"cd", -- 1230
         x"71",  x"00",  x"20",  x"7c",  x"e5",  x"c5",  x"13",  x"1a", -- 1238
         x"b7",  x"28",  x"09",  x"cd",  x"7f",  x"00",  x"28",  x"f6", -- 1240
         x"c1",  x"e1",  x"18",  x"e5",  x"c1",  x"d1",  x"ed",  x"5b", -- 1248
         x"1e",  x"00",  x"2b",  x"ed",  x"52",  x"c8",  x"44",  x"4d", -- 1250
         x"ed",  x"5b",  x"1c",  x"00",  x"2a",  x"1e",  x"00",  x"cd", -- 1258
         x"63",  x"00",  x"ed",  x"53",  x"1c",  x"00",  x"22",  x"1e", -- 1260
         x"00",  x"11",  x"01",  x"00",  x"e5",  x"cd",  x"9f",  x"d6", -- 1268
         x"e1",  x"ed",  x"5b",  x"1e",  x"00",  x"af",  x"ed",  x"52", -- 1270
         x"45",  x"4f",  x"28",  x"1e",  x"21",  x"24",  x"00",  x"be", -- 1278
         x"23",  x"28",  x"04",  x"10",  x"fa",  x"18",  x"13",  x"eb", -- 1280
         x"cd",  x"86",  x"00",  x"eb",  x"13",  x"0c",  x"fe",  x"09", -- 1288
         x"20",  x"06",  x"79",  x"c6",  x"07",  x"e6",  x"78",  x"4f", -- 1290
         x"10",  x"ed",  x"79",  x"fe",  x"50",  x"38",  x"02",  x"3e", -- 1298
         x"4f",  x"6f",  x"26",  x"00",  x"22",  x"20",  x"00",  x"3e", -- 12A0
         x"03",  x"bc",  x"c8",  x"11",  x"01",  x"00",  x"cd",  x"9f", -- 12A8
         x"d6",  x"c8",  x"2a",  x"20",  x"00",  x"24",  x"18",  x"ec", -- 12B0
         x"11",  x"00",  x"00",  x"cd",  x"4a",  x"d6",  x"21",  x"00", -- 12B8
         x"15",  x"22",  x"20",  x"00",  x"55",  x"5c",  x"cd",  x"9f", -- 12C0
         x"d6",  x"c9",  x"dd",  x"dd",  x"45",  x"44",  x"49",  x"54", -- 12C8
         x"1f",  x"cd",  x"9b",  x"de",  x"21",  x"9c",  x"cb",  x"e3", -- 12D0
         x"2a",  x"e7",  x"bf",  x"11",  x"dd",  x"dd",  x"a7",  x"ed", -- 12D8
         x"52",  x"28",  x"04",  x"dd",  x"cb",  x"08",  x"be",  x"cd", -- 12E0
         x"37",  x"ca",  x"cd",  x"83",  x"c8",  x"cd",  x"ec",  x"d3", -- 12E8
         x"cd",  x"ed",  x"d7",  x"cd",  x"39",  x"d9",  x"cd",  x"17", -- 12F0
         x"d5",  x"2a",  x"1c",  x"00",  x"22",  x"d8",  x"b4",  x"2a", -- 12F8
         x"1e",  x"00",  x"22",  x"da",  x"b4",  x"30",  x"55",  x"cd", -- 1300
         x"05",  x"d7",  x"38",  x"6c",  x"2a",  x"1a",  x"00",  x"ed", -- 1308
         x"5b",  x"1e",  x"00",  x"ed",  x"52",  x"44",  x"4d",  x"19", -- 1310
         x"ed",  x"5b",  x"1a",  x"00",  x"28",  x"25",  x"2b",  x"cd", -- 1318
         x"86",  x"00",  x"fe",  x"0a",  x"20",  x"08",  x"2b",  x"cd", -- 1320
         x"86",  x"00",  x"fe",  x"0d",  x"28",  x"e1",  x"23",  x"23", -- 1328
         x"ed",  x"5b",  x"1a",  x"00",  x"1b",  x"b7",  x"ed",  x"52", -- 1330
         x"30",  x"0d",  x"28",  x"0b",  x"19",  x"03",  x"03",  x"cd", -- 1338
         x"6a",  x"00",  x"13",  x"ed",  x"53",  x"1e",  x"00",  x"cd", -- 1340
         x"96",  x"ca",  x"21",  x"00",  x"ad",  x"11",  x"01",  x"ad", -- 1348
         x"01",  x"ff",  x"09",  x"36",  x"00",  x"ed",  x"b0",  x"dd", -- 1350
         x"cb",  x"08",  x"fe",  x"c9",  x"fe",  x"0d",  x"20",  x"02", -- 1358
         x"3e",  x"0e",  x"fe",  x"7f",  x"20",  x"02",  x"3e",  x"5f", -- 1360
         x"cd",  x"8d",  x"d3",  x"2a",  x"a0",  x"b7",  x"22",  x"20", -- 1368
         x"00",  x"3a",  x"22",  x"00",  x"b7",  x"ca",  x"f3",  x"d2", -- 1370
         x"cd",  x"fe",  x"d4",  x"cd",  x"40",  x"d8",  x"2a",  x"d8", -- 1378
         x"b4",  x"22",  x"1c",  x"00",  x"2a",  x"da",  x"b4",  x"22", -- 1380
         x"1e",  x"00",  x"c3",  x"f3",  x"d2",  x"fe",  x"20",  x"38", -- 1388
         x"33",  x"21",  x"3e",  x"00",  x"cb",  x"66",  x"20",  x"2c", -- 1390
         x"08",  x"cd",  x"c7",  x"d3",  x"d8",  x"08",  x"ed",  x"5b", -- 1398
         x"a0",  x"b7",  x"cd",  x"60",  x"c5",  x"46",  x"77",  x"cd", -- 13A0
         x"b4",  x"c5",  x"78",  x"a7",  x"28",  x"0e",  x"1c",  x"cd", -- 13A8
         x"60",  x"c5",  x"30",  x"f1",  x"1e",  x"00",  x"14",  x"cd", -- 13B0
         x"60",  x"c5",  x"30",  x"e9",  x"ed",  x"5b",  x"a0",  x"b7", -- 13B8
         x"cd",  x"60",  x"c5",  x"7e",  x"c3",  x"36",  x"c6",  x"0e", -- 13C0
         x"01",  x"c5",  x"ed",  x"5b",  x"a0",  x"b7",  x"cd",  x"60", -- 13C8
         x"c5",  x"eb",  x"21",  x"d0",  x"b4",  x"af",  x"ed",  x"52", -- 13D0
         x"44",  x"4d",  x"eb",  x"d1",  x"ed",  x"b1",  x"37",  x"c0", -- 13D8
         x"3f",  x"e2",  x"e8",  x"d3",  x"1d",  x"20",  x"f5",  x"c9", -- 13E0
         x"1d",  x"c8",  x"37",  x"c9",  x"ed",  x"5b",  x"18",  x"00", -- 13E8
         x"1b",  x"2a",  x"1c",  x"00",  x"a7",  x"ed",  x"52",  x"44", -- 13F0
         x"4d",  x"eb",  x"11",  x"00",  x"00",  x"3e",  x"0d",  x"cd", -- 13F8
         x"71",  x"00",  x"20",  x"04",  x"13",  x"ea",  x"ff",  x"d3", -- 1400
         x"ed",  x"53",  x"12",  x"00",  x"c9",  x"3e",  x"16",  x"92", -- 1408
         x"47",  x"c4",  x"a6",  x"c7",  x"ed",  x"5b",  x"9e",  x"b7", -- 1410
         x"15",  x"1e",  x"00",  x"cd",  x"60",  x"c5",  x"ed",  x"4b", -- 1418
         x"1e",  x"00",  x"cd",  x"88",  x"d7",  x"ed",  x"5b",  x"a0", -- 1420
         x"b7",  x"c3",  x"e4",  x"c6",  x"3a",  x"3e",  x"00",  x"e6", -- 1428
         x"10",  x"20",  x"1c",  x"7b",  x"2f",  x"e6",  x"07",  x"3c", -- 1430
         x"47",  x"4f",  x"c5",  x"cd",  x"c9",  x"d3",  x"c1",  x"ed", -- 1438
         x"5b",  x"a0",  x"b7",  x"d8",  x"c5",  x"3e",  x"20",  x"cd", -- 1440
         x"9e",  x"d3",  x"36",  x"00",  x"c1",  x"10",  x"f5",  x"cd", -- 1448
         x"95",  x"c6",  x"7b",  x"e6",  x"07",  x"20",  x"f8",  x"c9", -- 1450
         x"3a",  x"3e",  x"00",  x"e6",  x"10",  x"20",  x"60",  x"3a", -- 1458
         x"9f",  x"b7",  x"3d",  x"ba",  x"20",  x"08",  x"cd",  x"04", -- 1460
         x"c7",  x"15",  x"ed",  x"53",  x"a0",  x"b7",  x"2a",  x"1c", -- 1468
         x"00",  x"e5",  x"21",  x"80",  x"b4",  x"cd",  x"2b",  x"d7", -- 1470
         x"d1",  x"d4",  x"e8",  x"d6",  x"ed",  x"5b",  x"a0",  x"b7", -- 1478
         x"3a",  x"9f",  x"b7",  x"3d",  x"92",  x"3d",  x"47",  x"cd", -- 1480
         x"00",  x"c8",  x"ed",  x"5b",  x"a0",  x"b7",  x"2a",  x"10", -- 1488
         x"00",  x"62",  x"24",  x"7b",  x"bd",  x"30",  x"02",  x"2e", -- 1490
         x"00",  x"22",  x"a0",  x"b7",  x"45",  x"cd",  x"60",  x"c5", -- 1498
         x"4e",  x"af",  x"77",  x"cd",  x"b4",  x"c5",  x"d5",  x"14", -- 14A0
         x"58",  x"cd",  x"60",  x"c5",  x"79",  x"77",  x"cd",  x"b4", -- 14A8
         x"c5",  x"1c",  x"43",  x"d1",  x"1c",  x"7b",  x"fe",  x"51", -- 14B0
         x"20",  x"e3",  x"ed",  x"5b",  x"a0",  x"b7",  x"c9",  x"cd", -- 14B8
         x"d7",  x"c6",  x"3a",  x"10",  x"00",  x"5f",  x"c9",  x"11", -- 14C0
         x"00",  x"00",  x"cd",  x"60",  x"c5",  x"cd",  x"2b",  x"d7", -- 14C8
         x"3a",  x"a1",  x"b7",  x"3c",  x"32",  x"9f",  x"b7",  x"c3", -- 14D0
         x"87",  x"ce",  x"cd",  x"03",  x"f0",  x"0c",  x"d0",  x"fe", -- 14D8
         x"03",  x"37",  x"c8",  x"fe",  x"13",  x"37",  x"3f",  x"c0", -- 14E0
         x"cd",  x"17",  x"d5",  x"d8",  x"18",  x"f5",  x"2a",  x"a0", -- 14E8
         x"b7",  x"e5",  x"cd",  x"89",  x"ca",  x"af",  x"32",  x"a1", -- 14F0
         x"b7",  x"cd",  x"21",  x"d5",  x"18",  x"0e",  x"2a",  x"a0", -- 14F8
         x"b7",  x"e5",  x"cd",  x"89",  x"ca",  x"af",  x"32",  x"a1", -- 1500
         x"b7",  x"cd",  x"41",  x"d5",  x"cd",  x"17",  x"d5",  x"cd", -- 1508
         x"6e",  x"d9",  x"e1",  x"22",  x"a0",  x"b7",  x"c9",  x"cd", -- 1510
         x"03",  x"f0",  x"04",  x"fe",  x"03",  x"37",  x"c8",  x"3f", -- 1518
         x"c9",  x"cd",  x"03",  x"f0",  x"23",  x"0d",  x"09",  x"3e", -- 1520
         x"3e",  x"3e",  x"3e",  x"20",  x"42",  x"6c",  x"6f",  x"63", -- 1528
         x"6b",  x"2d",  x"4d",  x"61",  x"72",  x"6b",  x"65",  x"6e", -- 1530
         x"3f",  x"20",  x"3c",  x"3c",  x"3c",  x"3c",  x"08",  x"00", -- 1538
         x"c9",  x"cd",  x"03",  x"f0",  x"23",  x"0d",  x"09",  x"3e", -- 1540
         x"3e",  x"3e",  x"3e",  x"20",  x"53",  x"70",  x"65",  x"69", -- 1548
         x"63",  x"68",  x"65",  x"72",  x"20",  x"76",  x"6f",  x"6c", -- 1550
         x"6c",  x"20",  x"3c",  x"3c",  x"3c",  x"3c",  x"08",  x"00", -- 1558
         x"af",  x"32",  x"22",  x"00",  x"c9",  x"cd",  x"03",  x"f0", -- 1560
         x"23",  x"20",  x"28",  x"59",  x"2f",  x"4e",  x"29",  x"20", -- 1568
         x"3f",  x"20",  x"00",  x"cd",  x"17",  x"d5",  x"38",  x"0c", -- 1570
         x"cd",  x"4c",  x"db",  x"fe",  x"59",  x"28",  x"05",  x"fe", -- 1578
         x"4e",  x"20",  x"f0",  x"37",  x"f5",  x"cd",  x"8c",  x"ce", -- 1580
         x"cd",  x"87",  x"ce",  x"f1",  x"c9",  x"3a",  x"df",  x"b7", -- 1588
         x"f5",  x"af",  x"32",  x"df",  x"b7",  x"78",  x"32",  x"a0", -- 1590
         x"b7",  x"cd",  x"17",  x"d5",  x"30",  x"09",  x"cd",  x"87", -- 1598
         x"ce",  x"f1",  x"32",  x"df",  x"b7",  x"37",  x"c9",  x"fe", -- 15A0
         x"2e",  x"28",  x"23",  x"fe",  x"05",  x"28",  x"24",  x"fe", -- 15A8
         x"20",  x"30",  x"2a",  x"fe",  x"08",  x"28",  x"26",  x"fe", -- 15B0
         x"09",  x"28",  x"22",  x"fe",  x"0d",  x"20",  x"da",  x"3a", -- 15B8
         x"a1",  x"b7",  x"57",  x"58",  x"cd",  x"03",  x"f0",  x"32", -- 15C0
         x"f1",  x"32",  x"df",  x"b7",  x"a7",  x"c9",  x"79",  x"fe", -- 15C8
         x"10",  x"20",  x"08",  x"78",  x"c6",  x"08",  x"32",  x"a0", -- 15D0
         x"b7",  x"18",  x"06",  x"3e",  x"2e",  x"cd",  x"03",  x"f0", -- 15D8
         x"00",  x"21",  x"a0",  x"b7",  x"7e",  x"b8",  x"30",  x"01", -- 15E0
         x"78",  x"b9",  x"38",  x"01",  x"79",  x"77",  x"18",  x"a9", -- 15E8
         x"cd",  x"03",  x"f0",  x"23",  x"0a",  x"0b",  x"4e",  x"61", -- 15F0
         x"6d",  x"65",  x"20",  x"3a",  x"00",  x"21",  x"f5",  x"b7", -- 15F8
         x"06",  x"08",  x"cd",  x"2b",  x"d6",  x"7e",  x"fe",  x"21", -- 1600
         x"38",  x"07",  x"06",  x"03",  x"cd",  x"2b",  x"d6",  x"18", -- 1608
         x"08",  x"cd",  x"03",  x"f0",  x"23",  x"54",  x"58",  x"54", -- 1610
         x"00",  x"01",  x"10",  x"06",  x"cd",  x"8d",  x"d5",  x"d8", -- 1618
         x"11",  x"00",  x"00",  x"d5",  x"01",  x"0b",  x"00",  x"ed", -- 1620
         x"b0",  x"e1",  x"c9",  x"7e",  x"e6",  x"7f",  x"23",  x"cd", -- 1628
         x"03",  x"f0",  x"42",  x"10",  x"f6",  x"c9",  x"11",  x"80", -- 1630
         x"b7",  x"af",  x"1d",  x"12",  x"20",  x"fc",  x"dd",  x"73", -- 1638
         x"05",  x"dd",  x"72",  x"06",  x"01",  x"0b",  x"00",  x"ed", -- 1640
         x"b0",  x"c9",  x"2a",  x"1a",  x"00",  x"ed",  x"4b",  x"1e", -- 1648
         x"00",  x"af",  x"ed",  x"42",  x"44",  x"4d",  x"c8",  x"2a", -- 1650
         x"12",  x"00",  x"e5",  x"2a",  x"1e",  x"00",  x"3e",  x"0d", -- 1658
         x"cd",  x"71",  x"00",  x"20",  x"13",  x"1b",  x"e3",  x"23", -- 1660
         x"e3",  x"e2",  x"78",  x"d6",  x"7a",  x"b3",  x"20",  x"ee", -- 1668
         x"cd",  x"86",  x"00",  x"fe",  x"0a",  x"20",  x"01",  x"23", -- 1670
         x"cd",  x"80",  x"d6",  x"e1",  x"22",  x"12",  x"00",  x"c9", -- 1678
         x"ed",  x"5b",  x"1e",  x"00",  x"d5",  x"af",  x"ed",  x"52", -- 1680
         x"44",  x"4d",  x"e1",  x"ed",  x"5b",  x"1c",  x"00",  x"28", -- 1688
         x"03",  x"cd",  x"63",  x"00",  x"ed",  x"53",  x"1c",  x"00", -- 1690
         x"22",  x"1e",  x"00",  x"c9",  x"cd",  x"e2",  x"cd",  x"2a", -- 1698
         x"1c",  x"00",  x"ed",  x"4b",  x"18",  x"00",  x"af",  x"ed", -- 16A0
         x"42",  x"44",  x"4d",  x"c8",  x"03",  x"2a",  x"12",  x"00", -- 16A8
         x"e5",  x"2a",  x"1c",  x"00",  x"2b",  x"cd",  x"86",  x"00", -- 16B0
         x"fe",  x"0a",  x"20",  x"02",  x"2b",  x"0b",  x"cd",  x"86", -- 16B8
         x"00",  x"fe",  x"0d",  x"20",  x"02",  x"2b",  x"0b",  x"3e", -- 16C0
         x"0d",  x"cd",  x"78",  x"00",  x"1b",  x"e3",  x"2b",  x"e3", -- 16C8
         x"20",  x"08",  x"e2",  x"d9",  x"d6",  x"7a",  x"b3",  x"20", -- 16D0
         x"ee",  x"23",  x"23",  x"cd",  x"86",  x"00",  x"fe",  x"0a", -- 16D8
         x"20",  x"01",  x"23",  x"eb",  x"e1",  x"22",  x"12",  x"00", -- 16E0
         x"2a",  x"1c",  x"00",  x"e5",  x"af",  x"ed",  x"52",  x"44", -- 16E8
         x"4d",  x"e1",  x"ed",  x"5b",  x"1e",  x"00",  x"1b",  x"2b", -- 16F0
         x"c4",  x"6a",  x"00",  x"13",  x"ed",  x"53",  x"1e",  x"00", -- 16F8
         x"23",  x"22",  x"1c",  x"00",  x"c9",  x"2a",  x"1e",  x"00", -- 1700
         x"22",  x"da",  x"b4",  x"2a",  x"1c",  x"00",  x"22",  x"d8", -- 1708
         x"b4",  x"2a",  x"1c",  x"00",  x"e5",  x"11",  x"00",  x"00", -- 1710
         x"cd",  x"60",  x"c5",  x"06",  x"17",  x"c5",  x"cd",  x"2b", -- 1718
         x"d7",  x"c1",  x"38",  x"05",  x"10",  x"f7",  x"d1",  x"18", -- 1720
         x"bf",  x"d1",  x"c9",  x"ed",  x"5b",  x"1c",  x"00",  x"06", -- 1728
         x"50",  x"0e",  x"00",  x"7e",  x"23",  x"a7",  x"28",  x"0d", -- 1730
         x"cd",  x"73",  x"d7",  x"d8",  x"10",  x"f3",  x"18",  x"08", -- 1738
         x"7e",  x"23",  x"a7",  x"20",  x"14",  x"0c",  x"10",  x"f8", -- 1740
         x"3e",  x"0d",  x"cd",  x"73",  x"d7",  x"d8",  x"3e",  x"0a", -- 1748
         x"cd",  x"73",  x"d7",  x"d8",  x"ed",  x"53",  x"1c",  x"00", -- 1750
         x"c9",  x"f5",  x"79",  x"c6",  x"07",  x"cb",  x"3f",  x"cb", -- 1758
         x"3f",  x"cb",  x"3f",  x"4f",  x"3e",  x"09",  x"cd",  x"73", -- 1760
         x"d7",  x"38",  x"06",  x"0d",  x"20",  x"f8",  x"f1",  x"18", -- 1768
         x"c7",  x"c1",  x"c9",  x"e5",  x"2a",  x"1e",  x"00",  x"37", -- 1770
         x"ed",  x"52",  x"e1",  x"38",  x"07",  x"eb",  x"cd",  x"92", -- 1778
         x"00",  x"eb",  x"13",  x"c9",  x"32",  x"22",  x"00",  x"c9", -- 1780
         x"7b",  x"fe",  x"50",  x"30",  x"33",  x"cd",  x"8c",  x"00", -- 1788
         x"fe",  x"03",  x"28",  x"4e",  x"03",  x"fe",  x"20",  x"38", -- 1790
         x"07",  x"cd",  x"b1",  x"c5",  x"23",  x"1c",  x"18",  x"e8", -- 1798
         x"fe",  x"09",  x"20",  x"10",  x"cd",  x"b0",  x"c5",  x"23", -- 17A0
         x"1c",  x"7b",  x"fe",  x"50",  x"30",  x"12",  x"e6",  x"07", -- 17A8
         x"20",  x"f2",  x"18",  x"d4",  x"fe",  x"0d",  x"28",  x"1d", -- 17B0
         x"fe",  x"0a",  x"28",  x"0f",  x"fe",  x"03",  x"18",  x"d9", -- 17B8
         x"cd",  x"8c",  x"00",  x"fe",  x"0d",  x"28",  x"0e",  x"fe", -- 17C0
         x"0a",  x"20",  x"13",  x"03",  x"cd",  x"8c",  x"00",  x"fe", -- 17C8
         x"0d",  x"20",  x"0b",  x"18",  x"08",  x"03",  x"cd",  x"8c", -- 17D0
         x"00",  x"fe",  x"0a",  x"20",  x"01",  x"03",  x"ed",  x"43", -- 17D8
         x"1e",  x"00",  x"7b",  x"fe",  x"50",  x"d0",  x"cd",  x"b0", -- 17E0
         x"c5",  x"23",  x"1c",  x"18",  x"f5",  x"cd",  x"40",  x"d8", -- 17E8
         x"ed",  x"4b",  x"1e",  x"00",  x"11",  x"00",  x"00",  x"cd", -- 17F0
         x"60",  x"c5",  x"1e",  x"00",  x"cd",  x"88",  x"d7",  x"14", -- 17F8
         x"7a",  x"fe",  x"17",  x"20",  x"f5",  x"c3",  x"85",  x"c9", -- 1800
         x"00",  x"00",  x"ff",  x"00",  x"3f",  x"01",  x"ff",  x"00", -- 1808
         x"00",  x"00",  x"ed",  x"00",  x"3f",  x"01",  x"ed",  x"00", -- 1810
         x"00",  x"00",  x"ed",  x"00",  x"00",  x"00",  x"ff",  x"00", -- 1818
         x"3f",  x"01",  x"ee",  x"00",  x"3f",  x"01",  x"fe",  x"00", -- 1820
         x"6a",  x"00",  x"ee",  x"00",  x"6a",  x"00",  x"fe",  x"00", -- 1828
         x"aa",  x"00",  x"ee",  x"00",  x"aa",  x"00",  x"fe",  x"00", -- 1830
         x"ee",  x"00",  x"ee",  x"00",  x"ee",  x"00",  x"fe",  x"00", -- 1838
         x"cd",  x"89",  x"ca",  x"3e",  x"3c",  x"32",  x"d6",  x"b7", -- 1840
         x"21",  x"08",  x"d8",  x"06",  x"07",  x"c5",  x"11",  x"82", -- 1848
         x"b7",  x"01",  x"08",  x"00",  x"ed",  x"b0",  x"e5",  x"cd", -- 1850
         x"03",  x"f0",  x"3e",  x"e1",  x"c1",  x"10",  x"ee",  x"21", -- 1858
         x"01",  x"00",  x"22",  x"a0",  x"b7",  x"cd",  x"03",  x"f0", -- 1860
         x"23",  x"5a",  x"65",  x"69",  x"6c",  x"65",  x"3a",  x"20", -- 1868
         x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"53",  x"70", -- 1870
         x"61",  x"6c",  x"74",  x"65",  x"3a",  x"20",  x"00",  x"cd", -- 1878
         x"85",  x"d9",  x"3e",  x"1e",  x"32",  x"a0",  x"b7",  x"21", -- 1880
         x"3e",  x"00",  x"cb",  x"66",  x"20",  x"10",  x"cd",  x"03", -- 1888
         x"f0",  x"23",  x"45",  x"69",  x"6e",  x"66",  x"81",  x"67", -- 1890
         x"65",  x"6e",  x"20",  x"00",  x"18",  x"0e",  x"cd",  x"03", -- 1898
         x"f0",  x"23",  x"9a",  x"62",  x"65",  x"72",  x"73",  x"63", -- 18A0
         x"68",  x"72",  x"2e",  x"00",  x"3e",  x"2d",  x"32",  x"a0", -- 18A8
         x"b7",  x"cd",  x"03",  x"f0",  x"23",  x"5a",  x"53",  x"3a", -- 18B0
         x"00",  x"7e",  x"e6",  x"60",  x"20",  x"10",  x"cd",  x"03", -- 18B8
         x"f0",  x"23",  x"61",  x"6d",  x"65",  x"72",  x"69",  x"6b", -- 18C0
         x"61",  x"6e",  x"2e",  x"00",  x"18",  x"22",  x"d6",  x"20", -- 18C8
         x"20",  x"10",  x"cd",  x"03",  x"f0",  x"23",  x"64",  x"65", -- 18D0
         x"75",  x"74",  x"73",  x"63",  x"68",  x"20",  x"20",  x"00", -- 18D8
         x"18",  x"0e",  x"cd",  x"03",  x"f0",  x"23",  x"43",  x"41", -- 18E0
         x"4f",  x"53",  x"20",  x"20",  x"20",  x"20",  x"20",  x"00", -- 18E8
         x"3e",  x"40",  x"32",  x"a0",  x"b7",  x"21",  x"f5",  x"b7", -- 18F0
         x"06",  x"08",  x"cd",  x"2b",  x"d6",  x"3e",  x"2e",  x"cd", -- 18F8
         x"03",  x"f0",  x"00",  x"06",  x"03",  x"cd",  x"2b",  x"d6", -- 1900
         x"11",  x"28",  x"00",  x"dd",  x"cb",  x"08",  x"6e",  x"3e", -- 1908
         x"05",  x"20",  x"02",  x"3e",  x"20",  x"cd",  x"b4",  x"c5", -- 1910
         x"11",  x"00",  x"01",  x"2a",  x"10",  x"00",  x"06",  x"0a", -- 1918
         x"0e",  x"07",  x"7b",  x"bd",  x"20",  x"02",  x"0e",  x"02", -- 1920
         x"bc",  x"20",  x"02",  x"0e",  x"03",  x"79",  x"cd",  x"b4", -- 1928
         x"c5",  x"3e",  x"08",  x"83",  x"5f",  x"0e",  x"06",  x"10", -- 1930
         x"e9",  x"cd",  x"89",  x"ca",  x"21",  x"08",  x"00",  x"22", -- 1938
         x"a0",  x"b7",  x"2a",  x"21",  x"00",  x"26",  x"00",  x"ed", -- 1940
         x"5b",  x"12",  x"00",  x"19",  x"cd",  x"f6",  x"de",  x"cd", -- 1948
         x"03",  x"f0",  x"2b",  x"21",  x"16",  x"00",  x"22",  x"a0", -- 1950
         x"b7",  x"2a",  x"20",  x"00",  x"26",  x"00",  x"23",  x"cd", -- 1958
         x"f6",  x"de",  x"cd",  x"03",  x"f0",  x"2b",  x"ed",  x"5b", -- 1960
         x"20",  x"00",  x"ed",  x"53",  x"a0",  x"b7",  x"21",  x"00", -- 1968
         x"02",  x"22",  x"9c",  x"b7",  x"21",  x"50",  x"17",  x"22", -- 1970
         x"9e",  x"b7",  x"c9",  x"d5",  x"cd",  x"89",  x"ca",  x"cd", -- 1978
         x"85",  x"d9",  x"d1",  x"18",  x"e9",  x"dd",  x"cb",  x"08", -- 1980
         x"7e",  x"3e",  x"1d",  x"20",  x"02",  x"3e",  x"1f",  x"11", -- 1988
         x"1c",  x"00",  x"c3",  x"b4",  x"c5",  x"49",  x"4d",  x"50", -- 1990
         x"4f",  x"52",  x"54",  x"20",  x"20",  x"4b",  x"43",  x"43", -- 1998
         x"00",  x"dd",  x"dd",  x"49",  x"4d",  x"50",  x"4f",  x"52", -- 19A0
         x"54",  x"01",  x"21",  x"95",  x"d9",  x"cd",  x"03",  x"f0", -- 19A8
         x"23",  x"4c",  x"6f",  x"61",  x"64",  x"69",  x"6e",  x"67", -- 19B0
         x"20",  x"00",  x"e5",  x"cd",  x"03",  x"f0",  x"45",  x"cd", -- 19B8
         x"87",  x"ce",  x"e1",  x"11",  x"00",  x"00",  x"01",  x"0b", -- 19C0
         x"00",  x"ed",  x"b0",  x"21",  x"00",  x"00",  x"cd",  x"03", -- 19C8
         x"f0",  x"10",  x"d8",  x"c3",  x"00",  x"ba",  x"48",  x"49", -- 19D0
         x"4c",  x"46",  x"45",  x"20",  x"20",  x"20",  x"4b",  x"43", -- 19D8
         x"43",  x"00",  x"dd",  x"dd",  x"48",  x"45",  x"4c",  x"50", -- 19E0
         x"01",  x"21",  x"d6",  x"d9",  x"18",  x"bf",  x"eb",  x"b7", -- 19E8
         x"ed",  x"52",  x"4d",  x"44",  x"03",  x"eb",  x"3e",  x"1c", -- 19F0
         x"cd",  x"71",  x"00",  x"c0",  x"54",  x"5d",  x"3e",  x"1e", -- 19F8
         x"cd",  x"71",  x"00",  x"2b",  x"eb",  x"c9",  x"dd",  x"dd", -- 1A00
         x"50",  x"53",  x"41",  x"56",  x"45",  x"1f",  x"cd",  x"9c", -- 1A08
         x"d6",  x"2a",  x"1e",  x"00",  x"e5",  x"ed",  x"5b",  x"1a", -- 1A10
         x"00",  x"d5",  x"cd",  x"ee",  x"d9",  x"28",  x"0c",  x"d1", -- 1A18
         x"e1",  x"cd",  x"03",  x"f0",  x"20",  x"cd",  x"21",  x"d5", -- 1A20
         x"c3",  x"87",  x"ce",  x"22",  x"1e",  x"00",  x"ed",  x"53", -- 1A28
         x"1a",  x"00",  x"2a",  x"1a",  x"00",  x"cd",  x"86",  x"00", -- 1A30
         x"e5",  x"f5",  x"3e",  x"03",  x"cd",  x"92",  x"00",  x"cd", -- 1A38
         x"f4",  x"cd",  x"f1",  x"e1",  x"cd",  x"92",  x"00",  x"e1", -- 1A40
         x"22",  x"1a",  x"00",  x"e1",  x"22",  x"1e",  x"00",  x"c9", -- 1A48
         x"dd",  x"dd",  x"50",  x"50",  x"52",  x"49",  x"4e",  x"54", -- 1A50
         x"01",  x"cd",  x"e9",  x"d0",  x"d8",  x"cd",  x"9c",  x"d6", -- 1A58
         x"2a",  x"1e",  x"00",  x"e5",  x"ed",  x"5b",  x"1a",  x"00", -- 1A60
         x"d5",  x"cd",  x"ee",  x"d9",  x"20",  x"b1",  x"22",  x"1e", -- 1A68
         x"00",  x"ed",  x"53",  x"1a",  x"00",  x"2a",  x"1a",  x"00", -- 1A70
         x"cd",  x"86",  x"00",  x"e5",  x"f5",  x"3e",  x"03",  x"cd", -- 1A78
         x"92",  x"00",  x"cd",  x"0f",  x"d0",  x"18",  x"bb",  x"01", -- 1A80
         x"27",  x"06",  x"cd",  x"8d",  x"d5",  x"d8",  x"f5",  x"cd", -- 1A88
         x"87",  x"ce",  x"f1",  x"c9",  x"dd",  x"dd",  x"52",  x"45", -- 1A90
         x"50",  x"4c",  x"41",  x"43",  x"45",  x"01",  x"b7",  x"cc", -- 1A98
         x"9c",  x"d6",  x"cd",  x"03",  x"f0",  x"23",  x"0a",  x"0a", -- 1AA0
         x"0b",  x"0b",  x"46",  x"69",  x"6e",  x"64",  x"20",  x"3a", -- 1AA8
         x"00",  x"cd",  x"87",  x"da",  x"d8",  x"7e",  x"b7",  x"c8", -- 1AB0
         x"22",  x"14",  x"00",  x"cd",  x"03",  x"f0",  x"23",  x"52", -- 1AB8
         x"65",  x"70",  x"6c",  x"2e",  x"3a",  x"00",  x"cd",  x"87", -- 1AC0
         x"da",  x"d8",  x"22",  x"16",  x"00",  x"fd",  x"26",  x"00", -- 1AC8
         x"2a",  x"1a",  x"00",  x"ed",  x"5b",  x"1e",  x"00",  x"b7", -- 1AD0
         x"ed",  x"52",  x"c8",  x"44",  x"4d",  x"eb",  x"ed",  x"5b", -- 1AD8
         x"14",  x"00",  x"1a",  x"cd",  x"71",  x"00",  x"e2",  x"fe", -- 1AE0
         x"da",  x"c5",  x"e5",  x"13",  x"1a",  x"b7",  x"28",  x"2d", -- 1AE8
         x"cd",  x"7f",  x"00",  x"e2",  x"fc",  x"da",  x"28",  x"f3", -- 1AF0
         x"e1",  x"c1",  x"18",  x"e2",  x"e1",  x"c1",  x"11",  x"01", -- 1AF8
         x"00",  x"cd",  x"9f",  x"d6",  x"fd",  x"7c",  x"cd",  x"03", -- 1B00
         x"f0",  x"1c",  x"cd",  x"03",  x"f0",  x"23",  x"20",  x"52", -- 1B08
         x"65",  x"70",  x"6c",  x"61",  x"63",  x"65",  x"73",  x"0d", -- 1B10
         x"0b",  x"0b",  x"0b",  x"00",  x"c9",  x"e3",  x"2b",  x"c5", -- 1B18
         x"cd",  x"80",  x"d6",  x"ed",  x"5b",  x"1c",  x"00",  x"c1", -- 1B20
         x"e1",  x"e5",  x"22",  x"1e",  x"00",  x"2a",  x"16",  x"00", -- 1B28
         x"7e",  x"a7",  x"28",  x"09",  x"23",  x"eb",  x"cd",  x"92", -- 1B30
         x"00",  x"eb",  x"13",  x"18",  x"f3",  x"ed",  x"53",  x"1c", -- 1B38
         x"00",  x"fd",  x"7c",  x"c6",  x"01",  x"27",  x"fd",  x"67", -- 1B40
         x"e1",  x"d1",  x"18",  x"92",  x"fe",  x"41",  x"d8",  x"fe", -- 1B48
         x"5b",  x"3f",  x"d0",  x"fe",  x"61",  x"d8",  x"fe",  x"7b", -- 1B50
         x"3f",  x"d8",  x"e6",  x"df",  x"c9",  x"79",  x"cb",  x"3f", -- 1B58
         x"f6",  x"10",  x"21",  x"a2",  x"b7",  x"cb",  x"de",  x"e5", -- 1B60
         x"cd",  x"91",  x"d3",  x"e1",  x"cb",  x"9e",  x"ed",  x"5b", -- 1B68
         x"a0",  x"b7",  x"ed",  x"53",  x"20",  x"00",  x"c3",  x"39", -- 1B70
         x"d9",  x"3e",  x"0c",  x"21",  x"3e",  x"0e",  x"21",  x"3e", -- 1B78
         x"0f",  x"21",  x"3e",  x"1c",  x"21",  x"3e",  x"1d",  x"21", -- 1B80
         x"3e",  x"1e",  x"21",  x"3e",  x"1f",  x"18",  x"d3",  x"21", -- 1B88
         x"00",  x"00",  x"22",  x"9c",  x"b7",  x"22",  x"a0",  x"b7", -- 1B90
         x"cd",  x"03",  x"f0",  x"23",  x"5a",  x"65",  x"69",  x"63", -- 1B98
         x"68",  x"65",  x"6e",  x"20",  x"61",  x"75",  x"73",  x"77", -- 1BA0
         x"84",  x"68",  x"6c",  x"65",  x"6e",  x"20",  x"75",  x"6e", -- 1BA8
         x"64",  x"20",  x"42",  x"52",  x"4b",  x"2f",  x"45",  x"6e", -- 1BB0
         x"64",  x"65",  x"72",  x"3a",  x"00",  x"3e",  x"b0",  x"06", -- 1BB8
         x"30",  x"cd",  x"03",  x"f0",  x"00",  x"3c",  x"10",  x"f9", -- 1BC0
         x"3e",  x"80",  x"06",  x"30",  x"cd",  x"03",  x"f0",  x"00", -- 1BC8
         x"3c",  x"10",  x"f9",  x"3e",  x"e0",  x"06",  x"20",  x"cd", -- 1BD0
         x"03",  x"f0",  x"00",  x"3c",  x"10",  x"f9",  x"2a",  x"de", -- 1BD8
         x"b4",  x"22",  x"a0",  x"b7",  x"cd",  x"17",  x"d5",  x"38", -- 1BE0
         x"60",  x"2a",  x"a0",  x"b7",  x"fe",  x"08",  x"20",  x"14", -- 1BE8
         x"7c",  x"a7",  x"7d",  x"20",  x"07",  x"fe",  x"20",  x"28", -- 1BF0
         x"eb",  x"2d",  x"18",  x"e5",  x"a7",  x"20",  x"fa",  x"21", -- 1BF8
         x"4f",  x"00",  x"18",  x"dd",  x"fe",  x"09",  x"20",  x"15", -- 1C00
         x"7c",  x"a7",  x"7d",  x"28",  x"07",  x"fe",  x"4f",  x"28", -- 1C08
         x"d3",  x"2c",  x"18",  x"cd",  x"fe",  x"4f",  x"20",  x"f9", -- 1C10
         x"21",  x"00",  x"01",  x"18",  x"c4",  x"fe",  x"0a",  x"20", -- 1C18
         x"07",  x"7c",  x"3d",  x"28",  x"bf",  x"24",  x"18",  x"b9", -- 1C20
         x"fe",  x"0b",  x"20",  x"0c",  x"7c",  x"a7",  x"28",  x"b4", -- 1C28
         x"7d",  x"fe",  x"20",  x"38",  x"af",  x"25",  x"18",  x"a9", -- 1C30
         x"fe",  x"0d",  x"20",  x"a8",  x"eb",  x"cd",  x"60",  x"c5", -- 1C38
         x"7e",  x"f5",  x"cd",  x"49",  x"dc",  x"f1",  x"c3",  x"62", -- 1C40
         x"db",  x"2a",  x"a0",  x"b7",  x"22",  x"de",  x"b4",  x"3e", -- 1C48
         x"02",  x"32",  x"9f",  x"b7",  x"cd",  x"83",  x"c8",  x"c3", -- 1C50
         x"82",  x"c9",  x"21",  x"10",  x"00",  x"18",  x"03",  x"21", -- 1C58
         x"11",  x"00",  x"7b",  x"e6",  x"f8",  x"77",  x"18",  x"ef", -- 1C60
         x"cd",  x"84",  x"dc",  x"cd",  x"ec",  x"d3",  x"c3",  x"ed", -- 1C68
         x"d7",  x"cd",  x"4e",  x"dd",  x"18",  x"f5",  x"2a",  x"12", -- 1C70
         x"00",  x"22",  x"dc",  x"b4",  x"cd",  x"84",  x"dc",  x"d4", -- 1C78
         x"5a",  x"dd",  x"18",  x"e7",  x"cd",  x"60",  x"c5",  x"7e", -- 1C80
         x"32",  x"e0",  x"b4",  x"3e",  x"1a",  x"77",  x"cd",  x"05", -- 1C88
         x"d7",  x"30",  x"10",  x"ed",  x"5b",  x"20",  x"00",  x"cd", -- 1C90
         x"60",  x"c5",  x"3a",  x"e0",  x"b4",  x"77",  x"cd",  x"fe", -- 1C98
         x"d4",  x"37",  x"c9",  x"ed",  x"5b",  x"1e",  x"00",  x"2a", -- 1CA0
         x"1a",  x"00",  x"ed",  x"52",  x"44",  x"4d",  x"eb",  x"3e", -- 1CA8
         x"1a",  x"cd",  x"71",  x"00",  x"ed",  x"5b",  x"1e",  x"00", -- 1CB0
         x"ed",  x"52",  x"44",  x"4d",  x"0b",  x"eb",  x"ed",  x"5b", -- 1CB8
         x"1c",  x"00",  x"78",  x"b1",  x"c4",  x"63",  x"00",  x"ed", -- 1CC0
         x"53",  x"1c",  x"00",  x"3a",  x"e0",  x"b4",  x"cd",  x"92", -- 1CC8
         x"00",  x"a7",  x"20",  x"01",  x"23",  x"22",  x"1e",  x"00", -- 1CD0
         x"2a",  x"18",  x"00",  x"cd",  x"ee",  x"d9",  x"28",  x"14", -- 1CD8
         x"2a",  x"1e",  x"00",  x"ed",  x"5b",  x"1a",  x"00",  x"cd", -- 1CE0
         x"ee",  x"d9",  x"28",  x"08",  x"cd",  x"ee",  x"d4",  x"cd", -- 1CE8
         x"1b",  x"dd",  x"37",  x"c9",  x"d5",  x"eb",  x"ed",  x"52", -- 1CF0
         x"44",  x"4d",  x"2a",  x"1e",  x"00",  x"ed",  x"5b",  x"1c", -- 1CF8
         x"00",  x"ed",  x"52",  x"ed",  x"42",  x"e1",  x"30",  x"05", -- 1D00
         x"cd",  x"1b",  x"dd",  x"37",  x"c9",  x"2b",  x"ed",  x"5b", -- 1D08
         x"1e",  x"00",  x"1b",  x"cd",  x"6a",  x"00",  x"13",  x"ed", -- 1D10
         x"53",  x"1e",  x"00",  x"ed",  x"5b",  x"21",  x"00",  x"16", -- 1D18
         x"00",  x"3a",  x"20",  x"00",  x"a7",  x"28",  x"01",  x"1c", -- 1D20
         x"c3",  x"9f",  x"d6",  x"cd",  x"05",  x"d7",  x"30",  x"0b", -- 1D28
         x"cd",  x"fe",  x"d4",  x"cd",  x"40",  x"d8",  x"ed",  x"5b", -- 1D30
         x"20",  x"00",  x"c9",  x"cd",  x"b8",  x"d2",  x"cd",  x"ec", -- 1D38
         x"d3",  x"c3",  x"ed",  x"d7",  x"cd",  x"05",  x"d7",  x"38", -- 1D40
         x"e7",  x"cd",  x"9c",  x"d6",  x"18",  x"f0",  x"2a",  x"12", -- 1D48
         x"00",  x"22",  x"dc",  x"b4",  x"cd",  x"05",  x"d7",  x"da", -- 1D50
         x"fe",  x"d4",  x"11",  x"00",  x"00",  x"cd",  x"9f",  x"d6", -- 1D58
         x"2a",  x"1e",  x"00",  x"ed",  x"5b",  x"1a",  x"00",  x"cd", -- 1D60
         x"ee",  x"d9",  x"28",  x"05",  x"cd",  x"ee",  x"d4",  x"18", -- 1D68
         x"23",  x"d5",  x"ed",  x"5b",  x"1e",  x"00",  x"ed",  x"52", -- 1D70
         x"44",  x"4d",  x"eb",  x"ed",  x"5b",  x"18",  x"00",  x"78", -- 1D78
         x"b1",  x"c4",  x"63",  x"00",  x"1b",  x"ed",  x"53",  x"1c", -- 1D80
         x"00",  x"e1",  x"23",  x"22",  x"1e",  x"00",  x"11",  x"01", -- 1D88
         x"00",  x"cd",  x"9f",  x"d6",  x"cd",  x"ec",  x"d3",  x"2a", -- 1D90
         x"dc",  x"b4",  x"b7",  x"ed",  x"52",  x"c8",  x"38",  x"04", -- 1D98
         x"eb",  x"c3",  x"4a",  x"d6",  x"19",  x"eb",  x"b7",  x"ed", -- 1DA0
         x"52",  x"eb",  x"c3",  x"9f",  x"d6",  x"cd",  x"89",  x"ca", -- 1DA8
         x"af",  x"32",  x"a1",  x"b7",  x"32",  x"0d",  x"ad",  x"01", -- 1DB0
         x"0c",  x"08",  x"cd",  x"8d",  x"d5",  x"38",  x"41",  x"11", -- 1DB8
         x"08",  x"ad",  x"01",  x"00",  x"00",  x"1a",  x"e6",  x"df", -- 1DC0
         x"28",  x"1b",  x"1a",  x"fe",  x"30",  x"38",  x"e1",  x"fe", -- 1DC8
         x"3a",  x"30",  x"dd",  x"e6",  x"0f",  x"60",  x"69",  x"29", -- 1DD0
         x"29",  x"29",  x"09",  x"09",  x"06",  x"00",  x"4f",  x"09", -- 1DD8
         x"44",  x"4d",  x"13",  x"18",  x"e0",  x"2a",  x"12",  x"00", -- 1DE0
         x"11",  x"16",  x"00",  x"19",  x"ed",  x"42",  x"38",  x"13", -- 1DE8
         x"60",  x"69",  x"ed",  x"5b",  x"12",  x"00",  x"ed",  x"52", -- 1DF0
         x"38",  x"09",  x"65",  x"2e",  x"00",  x"22",  x"20",  x"00", -- 1DF8
         x"c3",  x"40",  x"d8",  x"ed",  x"43",  x"dc",  x"b4",  x"cd", -- 1E00
         x"6e",  x"d9",  x"cd",  x"05",  x"d7",  x"30",  x"11",  x"cd", -- 1E08
         x"fe",  x"d4",  x"2a",  x"d8",  x"b4",  x"22",  x"1c",  x"00", -- 1E10
         x"2a",  x"da",  x"b4",  x"22",  x"1e",  x"00",  x"18",  x"e0", -- 1E18
         x"cd",  x"94",  x"dd",  x"21",  x"00",  x"00",  x"22",  x"20", -- 1E20
         x"00",  x"c3",  x"ed",  x"d7",  x"cd",  x"89",  x"ca",  x"21", -- 1E28
         x"01",  x"00",  x"22",  x"a0",  x"b7",  x"cd",  x"03",  x"f0", -- 1E30
         x"23",  x"53",  x"75",  x"63",  x"68",  x"65",  x"3a",  x"00", -- 1E38
         x"11",  x"08",  x"00",  x"06",  x"11",  x"cd",  x"60",  x"c5", -- 1E40
         x"cd",  x"b0",  x"c5",  x"1c",  x"10",  x"f7",  x"01",  x"19", -- 1E48
         x"08",  x"cd",  x"8d",  x"d5",  x"38",  x"aa",  x"21",  x"08", -- 1E50
         x"ad",  x"11",  x"23",  x"00",  x"01",  x"1b",  x"00",  x"ed", -- 1E58
         x"b0",  x"cd",  x"40",  x"d8",  x"ed",  x"5b",  x"20",  x"00", -- 1E60
         x"3a",  x"23",  x"00",  x"b7",  x"c8",  x"cd",  x"05",  x"d7", -- 1E68
         x"38",  x"9d",  x"11",  x"01",  x"00",  x"cd",  x"4a",  x"d6", -- 1E70
         x"cd",  x"14",  x"d2",  x"cd",  x"ec",  x"d3",  x"cd",  x"ed", -- 1E78
         x"d7",  x"c3",  x"85",  x"c9",  x"ed",  x"5b",  x"a0",  x"b7", -- 1E80
         x"21",  x"48",  x"15",  x"22",  x"a0",  x"b7",  x"dd",  x"7e", -- 1E88
         x"01",  x"f6",  x"05",  x"dd",  x"77",  x"01",  x"d3",  x"84", -- 1E90
         x"cd",  x"17",  x"d5",  x"dd",  x"7e",  x"01",  x"e6",  x"fa", -- 1E98
         x"dd",  x"77",  x"01",  x"d3",  x"84",  x"ed",  x"53",  x"a0", -- 1EA0
         x"b7",  x"c9",  x"dd",  x"dd",  x"44",  x"49",  x"52",  x"1f", -- 1EA8
         x"cd",  x"21",  x"f0",  x"08",  x"c9",  x"dd",  x"dd",  x"43", -- 1EB0
         x"44",  x"1f",  x"cd",  x"21",  x"f0",  x"09",  x"c9",  x"dd", -- 1EB8
         x"dd",  x"52",  x"45",  x"4e",  x"1f",  x"cd",  x"21",  x"f0", -- 1EC0
         x"0b",  x"c9",  x"dd",  x"dd",  x"45",  x"52",  x"41",  x"1f", -- 1EC8
         x"cd",  x"21",  x"f0",  x"0a",  x"c9",  x"dd",  x"dd",  x"44", -- 1ED0
         x"45",  x"56",  x"49",  x"43",  x"45",  x"01",  x"a7",  x"28", -- 1ED8
         x"0e",  x"7d",  x"fe",  x"08",  x"30",  x"04",  x"cd",  x"f1", -- 1EE0
         x"de",  x"d0",  x"cd",  x"03",  x"f0",  x"19",  x"c9",  x"3e", -- 1EE8
         x"ff",  x"cd",  x"03",  x"f0",  x"49",  x"c9",  x"d5",  x"01", -- 1EF0
         x"f6",  x"ff",  x"11",  x"ff",  x"ff",  x"09",  x"13",  x"38", -- 1EF8
         x"fc",  x"01",  x"0a",  x"00",  x"09",  x"eb",  x"7c",  x"b5", -- 1F00
         x"c4",  x"f6",  x"de",  x"7b",  x"c6",  x"30",  x"cd",  x"03", -- 1F08
         x"f0",  x"00",  x"d1",  x"c9",  x"70",  x"c6",  x"8e",  x"c9", -- 1F10
         x"0d",  x"d4",  x"70",  x"c6",  x"70",  x"c6",  x"2c",  x"d4", -- 1F18
         x"68",  x"de",  x"70",  x"c6",  x"d1",  x"c8",  x"95",  x"c6", -- 1F20
         x"d7",  x"c6",  x"36",  x"c7",  x"ca",  x"c8",  x"c7",  x"c8", -- 1F28
         x"58",  x"d4",  x"1f",  x"c9",  x"c5",  x"c8",  x"68",  x"c8", -- 1F30
         x"45",  x"c8",  x"31",  x"c9",  x"7a",  x"c9",  x"70",  x"c6", -- 1F38
         x"7b",  x"d9",  x"70",  x"c6",  x"c2",  x"c6",  x"fb",  x"c8", -- 1F40
         x"70",  x"c9",  x"70",  x"c6",  x"70",  x"c6",  x"70",  x"c6", -- 1F48
         x"70",  x"c6",  x"c4",  x"c9",  x"82",  x"db",  x"2b",  x"dd", -- 1F50
         x"68",  x"dc",  x"8b",  x"db",  x"88",  x"db",  x"2c",  x"de", -- 1F58
         x"8f",  x"db",  x"84",  x"de",  x"70",  x"c6",  x"79",  x"db", -- 1F60
         x"71",  x"dc",  x"5a",  x"dc",  x"70",  x"c6",  x"7c",  x"db", -- 1F68
         x"70",  x"c6",  x"70",  x"c6",  x"70",  x"c6",  x"5f",  x"dc", -- 1F70
         x"70",  x"c6",  x"44",  x"dd",  x"85",  x"db",  x"76",  x"dc", -- 1F78
         x"70",  x"c6",  x"7f",  x"db",  x"70",  x"c6",  x"ad",  x"dd", -- 1F80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1F98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 1FF8
         x"6a",  x"3a",  x"39",  x"06",  x"66",  x"35",  x"ff",  x"00", -- 2000
         x"10",  x"22",  x"32",  x"27",  x"37",  x"08",  x"18",  x"2a", -- 2008
         x"3a",  x"2f",  x"3f",  x"76",  x"c3",  x"d3",  x"e3",  x"f3", -- 2010
         x"c9",  x"d9",  x"e9",  x"f9",  x"db",  x"eb",  x"fb",  x"cd", -- 2018
         x"ff",  x"cf",  x"01",  x"02",  x"03",  x"09",  x"0a",  x"0b", -- 2020
         x"c1",  x"c5",  x"ff",  x"c7",  x"00",  x"04",  x"05",  x"06", -- 2028
         x"c0",  x"c2",  x"c4",  x"c6",  x"ff",  x"c0",  x"00",  x"40", -- 2030
         x"80",  x"c0",  x"ff",  x"70",  x"71",  x"47",  x"57",  x"67", -- 2038
         x"4d",  x"4f",  x"5f",  x"6f",  x"ff",  x"cf",  x"42",  x"43", -- 2040
         x"4a",  x"4b",  x"ff",  x"c7",  x"40",  x"41",  x"44",  x"45", -- 2048
         x"ff",  x"e7",  x"a0",  x"a1",  x"a2",  x"ff",  x"f7",  x"b3", -- 2050
         x"a3",  x"ff",  x"d7",  x"46",  x"ff",  x"df",  x"56",  x"5e", -- 2058
         x"ff",  x"00",  x"00",  x"d8",  x"6a",  x"de",  x"51",  x"60", -- 2060
         x"da",  x"5b",  x"5c",  x"db",  x"61",  x"7a",  x"d5",  x"5a", -- 2068
         x"69",  x"98",  x"69",  x"b4",  x"26",  x"35",  x"b4",  x"1f", -- 2070
         x"35",  x"9f",  x"38",  x"b8",  x"1f",  x"cd",  x"38",  x"b8", -- 2078
         x"4d",  x"a8",  x"38",  x"29",  x"cd",  x"50",  x"6a",  x"cd", -- 2080
         x"50",  x"69",  x"df",  x"61",  x"68",  x"df",  x"4e",  x"69", -- 2088
         x"cd",  x"5a",  x"6a",  x"e4",  x"13",  x"db",  x"78",  x"cf", -- 2090
         x"76",  x"96",  x"ce",  x"4f",  x"98",  x"d0",  x"51",  x"9a", -- 2098
         x"d4",  x"58",  x"cd",  x"52",  x"df",  x"5c",  x"de",  x"58", -- 20A0
         x"4f",  x"de",  x"5e",  x"4f",  x"de",  x"58",  x"de",  x"5e", -- 20A8
         x"df",  x"58",  x"4d",  x"df",  x"5e",  x"4d",  x"df",  x"58", -- 20B0
         x"5f",  x"df",  x"5e",  x"58",  x"ce",  x"cf",  x"d0",  x"d1", -- 20B8
         x"d4",  x"d8",  x"d9",  x"cd",  x"da",  x"66",  x"e6",  x"da", -- 20C0
         x"4f",  x"cf",  x"dc",  x"5b",  x"dc",  x"51",  x"dc",  x"d9", -- 20C8
         x"d5",  x"d0",  x"d5",  x"5e",  x"d0",  x"5e",  x"b4",  x"1a", -- 20D0
         x"25",  x"35",  x"82",  x"d0",  x"56",  x"5a",  x"66",  x"2c", -- 20D8
         x"27",  x"80",  x"06",  x"09",  x"80",  x"06",  x"0b",  x"d0", -- 20E0
         x"4d",  x"4d",  x"df",  x"4f",  x"52",  x"d1",  x"7e",  x"1b", -- 20E8
         x"d6",  x"78",  x"27",  x"80",  x"08",  x"06",  x"80",  x"0a", -- 20F0
         x"06",  x"cf",  x"5c",  x"58",  x"cf",  x"4f",  x"52",  x"d4", -- 20F8
         x"4d",  x"58",  x"60",  x"d6",  x"76",  x"26",  x"83",  x"25", -- 2100
         x"d1",  x"7e",  x"34",  x"1c",  x"35",  x"09",  x"d0",  x"55", -- 2108
         x"81",  x"d1",  x"64",  x"64",  x"d6",  x"76",  x"07",  x"80", -- 2110
         x"08",  x"1a",  x"d5",  x"74",  x"0a",  x"25",  x"d1",  x"7e", -- 2118
         x"18",  x"38",  x"54",  x"58",  x"d1",  x"55",  x"cf",  x"4d", -- 2120
         x"58",  x"72",  x"26",  x"80",  x"08",  x"26",  x"80",  x"07", -- 2128
         x"0b",  x"84",  x"1f",  x"8d",  x"1a",  x"09",  x"80",  x"0a", -- 2130
         x"07",  x"85",  x"1f",  x"dc",  x"5b",  x"76",  x"1e",  x"dc", -- 2138
         x"61",  x"5f",  x"6e",  x"1e",  x"d6",  x"78",  x"23",  x"38", -- 2140
         x"27",  x"84",  x"21",  x"85",  x"21",  x"80",  x"21",  x"38", -- 2148
         x"25",  x"81",  x"2c",  x"22",  x"d6",  x"76",  x"22",  x"38", -- 2150
         x"26",  x"cf",  x"4d",  x"58",  x"72",  x"22",  x"38",  x"26", -- 2158
         x"9d",  x"25",  x"a0",  x"4d",  x"80",  x"21",  x"38",  x"29", -- 2160
         x"9d",  x"29",  x"de",  x"5f",  x"7a",  x"2b",  x"a0",  x"2c", -- 2168
         x"29",  x"2a",  x"ce",  x"55",  x"7a",  x"0c",  x"de",  x"51", -- 2170
         x"79",  x"0c",  x"2a",  x"df",  x"51",  x"7a",  x"0c",  x"2a", -- 2178
         x"d5",  x"5a",  x"52",  x"db",  x"60",  x"4f",  x"58",  x"80", -- 2180
         x"55",  x"0b",  x"80",  x"0a",  x"55",  x"de",  x"5e",  x"50", -- 2188
         x"81",  x"55",  x"80",  x"5e",  x"0b",  x"80",  x"0a",  x"5e", -- 2190
         x"de",  x"00",  x"90",  x"1a",  x"09",  x"80",  x"06",  x"09", -- 2198
         x"8e",  x"1a",  x"09",  x"80",  x"08",  x"06",  x"d5",  x"74", -- 21A0
         x"21",  x"38",  x"34",  x"4f",  x"35",  x"83",  x"34",  x"4f", -- 21A8
         x"35",  x"38",  x"21",  x"da",  x"51",  x"53",  x"81",  x"5a", -- 21B0
         x"d8",  x"50",  x"24",  x"cf",  x"5c",  x"24",  x"d5",  x"5a", -- 21B8
         x"24",  x"db",  x"60",  x"24",  x"db",  x"61",  x"60",  x"24", -- 21C0
         x"d5",  x"73",  x"3c",  x"d5",  x"73",  x"3d",  x"d5",  x"73", -- 21C8
         x"3e",  x"82",  x"d0",  x"68",  x"25",  x"d0",  x"68",  x"33", -- 21D0
         x"d0",  x"7d",  x"fe",  x"cb",  x"21",  x"01",  x"60",  x"20", -- 21D8
         x"1e",  x"2c",  x"cb",  x"49",  x"28",  x"20",  x"cb",  x"f9", -- 21E0
         x"13",  x"18",  x"1b",  x"0e",  x"00",  x"1a",  x"fe",  x"dd", -- 21E8
         x"20",  x"04",  x"0e",  x"02",  x"18",  x"06",  x"fe",  x"fd", -- 21F0
         x"20",  x"e0",  x"0e",  x"03",  x"13",  x"18",  x"ee",  x"fe", -- 21F8
         x"ed",  x"20",  x"04",  x"2d",  x"0e",  x"00",  x"13",  x"29", -- 2200
         x"46",  x"23",  x"6e",  x"1a",  x"a6",  x"23",  x"fd",  x"6f", -- 2208
         x"7e",  x"23",  x"fe",  x"ff",  x"28",  x"f5",  x"04",  x"fd", -- 2210
         x"bd",  x"20",  x"f5",  x"c5",  x"1a",  x"13",  x"fd",  x"6f", -- 2218
         x"0f",  x"0f",  x"0f",  x"e6",  x"07",  x"47",  x"f1",  x"18", -- 2220
         x"7a",  x"1a",  x"13",  x"6f",  x"26",  x"00",  x"fe",  x"80", -- 2228
         x"38",  x"01",  x"25",  x"19",  x"cd",  x"7e",  x"c3",  x"c3", -- 2230
         x"28",  x"c3",  x"1a",  x"13",  x"6f",  x"1a",  x"13",  x"67", -- 2238
         x"18",  x"f5",  x"1a",  x"13",  x"6f",  x"26",  x"00",  x"18", -- 2240
         x"ee",  x"07",  x"07",  x"07",  x"6f",  x"26",  x"00",  x"18", -- 2248
         x"e6",  x"c6",  x"3c",  x"fe",  x"2c",  x"38",  x"29",  x"d6", -- 2250
         x"0c",  x"fe",  x"20",  x"28",  x"10",  x"fe",  x"29",  x"20", -- 2258
         x"02",  x"cb",  x"91",  x"fe",  x"5b",  x"da",  x"0b",  x"cb", -- 2260
         x"d6",  x"1a",  x"cd",  x"0b",  x"cb",  x"cd",  x"00",  x"cb", -- 2268
         x"3a",  x"91",  x"b7",  x"a7",  x"c8",  x"3a",  x"a0",  x"b7", -- 2270
         x"fe",  x"0a",  x"d0",  x"cd",  x"00",  x"cb",  x"18",  x"f5", -- 2278
         x"e5",  x"21",  x"e4",  x"c2",  x"e5",  x"fe",  x"1d",  x"38", -- 2280
         x"1a",  x"fe",  x"25",  x"30",  x"2a",  x"fe",  x"1f",  x"38", -- 2288
         x"0c",  x"20",  x"02",  x"cb",  x"c0",  x"3d",  x"fe",  x"22", -- 2290
         x"38",  x"03",  x"cb",  x"90",  x"3d",  x"87",  x"87",  x"87", -- 2298
         x"d6",  x"db",  x"80",  x"cb",  x"49",  x"28",  x"54",  x"fe", -- 22A0
         x"1a",  x"20",  x"3b",  x"3e",  x"55",  x"cd",  x"53",  x"c2", -- 22A8
         x"79",  x"e6",  x"01",  x"c6",  x"64",  x"18",  x"9c",  x"c6", -- 22B0
         x"b8",  x"6f",  x"6e",  x"78",  x"cb",  x"79",  x"e9",  x"20", -- 22B8
         x"29",  x"fd",  x"7d",  x"e6",  x"07",  x"47",  x"3e",  x"20", -- 22C0
         x"18",  x"d3",  x"c8",  x"fd",  x"7d",  x"e6",  x"07",  x"fe", -- 22C8
         x"06",  x"20",  x"03",  x"cb",  x"71",  x"c0",  x"3e",  x"38", -- 22D0
         x"cd",  x"53",  x"c2",  x"18",  x"e4",  x"42",  x"3a",  x"29", -- 22D8
         x"51",  x"bf",  x"ca",  x"49",  x"e1",  x"c9",  x"fe",  x"2b", -- 22E0
         x"20",  x"11",  x"cb",  x"f1",  x"cb",  x"d1",  x"3e",  x"39", -- 22E8
         x"cb",  x"79",  x"28",  x"07",  x"1b",  x"1b",  x"cd",  x"fb", -- 22F0
         x"c2",  x"13",  x"c9",  x"3c",  x"21",  x"62",  x"c0",  x"23", -- 22F8
         x"cb",  x"7e",  x"28",  x"fb",  x"3d",  x"20",  x"f8",  x"7e", -- 2300
         x"e6",  x"7f",  x"cd",  x"53",  x"c2",  x"23",  x"cb",  x"7e", -- 2308
         x"28",  x"f5",  x"7d",  x"3d",  x"e6",  x"fe",  x"fe",  x"c0", -- 2310
         x"c0",  x"cb",  x"49",  x"c8",  x"cb",  x"71",  x"c0",  x"fd", -- 2318
         x"7d",  x"e6",  x"c7",  x"fe",  x"46",  x"c8",  x"18",  x"88", -- 2320
         x"cb",  x"51",  x"28",  x"12",  x"7d",  x"a7",  x"c8",  x"f2", -- 2328
         x"39",  x"c3",  x"ed",  x"44",  x"6f",  x"3e",  x"2d",  x"18", -- 2330
         x"02",  x"3e",  x"2b",  x"cd",  x"0b",  x"cb",  x"c5",  x"22", -- 2338
         x"97",  x"b7",  x"01",  x"40",  x"04",  x"21",  x"97",  x"b7", -- 2340
         x"af",  x"ed",  x"6f",  x"23",  x"ed",  x"6f",  x"a7",  x"20", -- 2348
         x"07",  x"cb",  x"71",  x"28",  x"03",  x"10",  x"ee",  x"04", -- 2350
         x"c6",  x"30",  x"fe",  x"3a",  x"38",  x"0e",  x"c6",  x"07", -- 2358
         x"cb",  x"71",  x"28",  x"08",  x"f5",  x"3e",  x"30",  x"cd", -- 2360
         x"0b",  x"cb",  x"0c",  x"f1",  x"cd",  x"0b",  x"cb",  x"0c", -- 2368
         x"cb",  x"b1",  x"10",  x"d1",  x"79",  x"e6",  x"fe",  x"c1", -- 2370
         x"c8",  x"3e",  x"48",  x"c3",  x"0b",  x"cb",  x"d5",  x"ed", -- 2378
         x"5b",  x"f5",  x"b7",  x"19",  x"d1",  x"c9",  x"7f",  x"dd", -- 2380
         x"fd",  x"a1",  x"3d",  x"3e",  x"3e",  x"02",  x"cd",  x"0b", -- 2388
         x"cb",  x"d5",  x"e1",  x"cd",  x"7e",  x"c3",  x"cd",  x"24", -- 2390
         x"cb",  x"cd",  x"00",  x"cb",  x"d5",  x"e1",  x"3a",  x"f4", -- 2398
         x"b7",  x"a7",  x"20",  x"69",  x"cd",  x"d9",  x"cd",  x"3a", -- 23A0
         x"f2",  x"b7",  x"cb",  x"5f",  x"28",  x"0f",  x"3e",  x"03", -- 23A8
         x"32",  x"f4",  x"b7",  x"0e",  x"00",  x"3e",  x"87",  x"cd", -- 23B0
         x"fb",  x"c2",  x"c3",  x"3a",  x"c2",  x"06",  x"00",  x"7e", -- 23B8
         x"fe",  x"cd",  x"20",  x"1a",  x"23",  x"7e",  x"fe",  x"21", -- 23C0
         x"28",  x"04",  x"fe",  x"03",  x"20",  x"17",  x"23",  x"7e", -- 23C8
         x"fe",  x"f0",  x"20",  x"1f",  x"23",  x"7e",  x"fe",  x"23", -- 23D0
         x"06",  x"04",  x"28",  x"02",  x"06",  x"01",  x"78",  x"32", -- 23D8
         x"f4",  x"b7",  x"c3",  x"eb",  x"c1",  x"fe",  x"0f",  x"20", -- 23E0
         x"0b",  x"23",  x"7e",  x"fe",  x"f0",  x"20",  x"04",  x"06", -- 23E8
         x"05",  x"18",  x"eb",  x"2b",  x"d5",  x"e5",  x"2a",  x"b0", -- 23F0
         x"b7",  x"11",  x"46",  x"00",  x"19",  x"d1",  x"1a",  x"be", -- 23F8
         x"20",  x"08",  x"23",  x"13",  x"1a",  x"be",  x"20",  x"02", -- 2400
         x"06",  x"02",  x"d1",  x"18",  x"d1",  x"d6",  x"02",  x"38", -- 2408
         x"32",  x"28",  x"0c",  x"32",  x"f4",  x"b7",  x"3d",  x"28", -- 2410
         x"06",  x"3d",  x"28",  x"2b",  x"af",  x"18",  x"36",  x"1a", -- 2418
         x"fe",  x"20",  x"38",  x"23",  x"fe",  x"80",  x"30",  x"1f", -- 2420
         x"3e",  x"86",  x"cd",  x"fb",  x"c2",  x"06",  x"14",  x"1a", -- 2428
         x"fe",  x"20",  x"38",  x"0a",  x"fe",  x"80",  x"30",  x"06", -- 2430
         x"cd",  x"0b",  x"cb",  x"13",  x"10",  x"f1",  x"3e",  x"27", -- 2438
         x"c3",  x"0b",  x"cb",  x"3c",  x"32",  x"f4",  x"b7",  x"1a", -- 2440
         x"a7",  x"20",  x"03",  x"32",  x"f4",  x"b7",  x"3e",  x"85", -- 2448
         x"0e",  x"00",  x"c3",  x"fb",  x"c2",  x"3e",  x"87",  x"0e", -- 2450
         x"00",  x"cd",  x"fb",  x"c2",  x"1a",  x"6f",  x"13",  x"1a", -- 2458
         x"67",  x"13",  x"19",  x"cd",  x"7e",  x"c3",  x"cd",  x"28", -- 2460
         x"c3",  x"21",  x"7b",  x"c4",  x"01",  x"00",  x"04",  x"7e", -- 2468
         x"23",  x"cd",  x"0b",  x"cb",  x"10",  x"f9",  x"af",  x"32", -- 2470
         x"f4",  x"b7",  x"c9",  x"2d",  x"24",  x"2d",  x"32",  x"7f", -- 2478
         x"7f",  x"44",  x"49",  x"53",  x"41",  x"53",  x"53",  x"01", -- 2480
         x"e5",  x"21",  x"f3",  x"db",  x"e3",  x"b7",  x"20",  x"2e", -- 2488
         x"cd",  x"03",  x"f0",  x"23",  x"0b",  x"09",  x"44",  x"49", -- 2490
         x"53",  x"41",  x"53",  x"53",  x"20",  x"41",  x"61",  x"64", -- 2498
         x"72",  x"20",  x"28",  x"5a",  x"65",  x"69",  x"6c",  x"65", -- 24A0
         x"6e",  x"20",  x"28",  x"41",  x"75",  x"73",  x"61",  x"64", -- 24A8
         x"72",  x"20",  x"28",  x"50",  x"72",  x"6f",  x"6c",  x"29", -- 24B0
         x"29",  x"29",  x"0d",  x"0a",  x"00",  x"c9",  x"c5",  x"4b", -- 24B8
         x"d1",  x"e5",  x"f5",  x"fe",  x"02",  x"38",  x"04",  x"79", -- 24C0
         x"b7",  x"20",  x"05",  x"ed",  x"4b",  x"9f",  x"b7",  x"0d", -- 24C8
         x"fd",  x"61",  x"f1",  x"fe",  x"03",  x"30",  x"02",  x"d1", -- 24D0
         x"d5",  x"e1",  x"eb",  x"b7",  x"ed",  x"52",  x"22",  x"f5", -- 24D8
         x"b7",  x"d5",  x"21",  x"86",  x"c3",  x"11",  x"f7",  x"b7", -- 24E0
         x"01",  x"06",  x"00",  x"ed",  x"b0",  x"fe",  x"04",  x"38", -- 24E8
         x"06",  x"2a",  x"88",  x"b7",  x"22",  x"fb",  x"b7",  x"d1", -- 24F0
         x"ed",  x"43",  x"f3",  x"b7",  x"3e",  x"09",  x"32",  x"91", -- 24F8
         x"b7",  x"fd",  x"44",  x"c5",  x"d5",  x"cd",  x"8c",  x"c3", -- 2500
         x"e1",  x"d5",  x"eb",  x"b7",  x"ed",  x"52",  x"7d",  x"fe", -- 2508
         x"04",  x"38",  x"02",  x"3e",  x"04",  x"4f",  x"3a",  x"a0", -- 2510
         x"b7",  x"fe",  x"19",  x"28",  x"12",  x"30",  x"1b",  x"3e", -- 2518
         x"09",  x"cd",  x"13",  x"cb",  x"18",  x"f0",  x"3e",  x"01", -- 2520
         x"32",  x"f4",  x"b7",  x"06",  x"01",  x"18",  x"d4",  x"41", -- 2528
         x"d5",  x"1a",  x"13",  x"cd",  x"03",  x"f0",  x"42",  x"10", -- 2530
         x"f8",  x"d1",  x"3a",  x"a0",  x"b7",  x"fe",  x"1e",  x"28", -- 2538
         x"09",  x"30",  x"0f",  x"3e",  x"09",  x"cd",  x"13",  x"cb", -- 2540
         x"18",  x"f0",  x"41",  x"1a",  x"13",  x"cd",  x"2f",  x"cb", -- 2548
         x"10",  x"f9",  x"d1",  x"cd",  x"57",  x"d2",  x"c1",  x"cd", -- 2550
         x"03",  x"f0",  x"2a",  x"d8",  x"10",  x"a5",  x"cd",  x"03", -- 2558
         x"f0",  x"04",  x"fe",  x"03",  x"c8",  x"fe",  x"0d",  x"28", -- 2560
         x"98",  x"fe",  x"0a",  x"28",  x"3b",  x"fe",  x"09",  x"28", -- 2568
         x"ba",  x"fe",  x"44",  x"28",  x"b1",  x"fe",  x"08",  x"28", -- 2570
         x"36",  x"fe",  x"0b",  x"20",  x"e1",  x"3a",  x"9f",  x"b7", -- 2578
         x"3d",  x"87",  x"47",  x"fd",  x"e5",  x"d5",  x"fd",  x"e1", -- 2580
         x"c5",  x"fd",  x"e5",  x"d1",  x"21",  x"f0",  x"ff",  x"19", -- 2588
         x"cd",  x"d9",  x"cd",  x"e5",  x"fd",  x"e1",  x"09",  x"af", -- 2590
         x"ed",  x"52",  x"19",  x"38",  x"f3",  x"c1",  x"10",  x"e8", -- 2598
         x"fd",  x"e5",  x"d1",  x"fd",  x"e1",  x"32",  x"f4",  x"b7", -- 25A0
         x"cd",  x"03",  x"f0",  x"2d",  x"c3",  x"01",  x"c5",  x"3a", -- 25A8
         x"9f",  x"b7",  x"18",  x"ce",  x"7f",  x"7f",  x"51",  x"4d", -- 25B0
         x"52",  x"01",  x"e5",  x"21",  x"f3",  x"db",  x"e3",  x"cd", -- 25B8
         x"03",  x"f0",  x"23",  x"02",  x"52",  x"65",  x"61",  x"73", -- 25C0
         x"73",  x"2e",  x"42",  x"65",  x"72",  x"65",  x"69",  x"63", -- 25C8
         x"68",  x"3a",  x"20",  x"00",  x"01",  x"1c",  x"0f",  x"cd", -- 25D0
         x"3d",  x"cf",  x"d8",  x"cd",  x"03",  x"f0",  x"18",  x"38", -- 25D8
         x"de",  x"2a",  x"97",  x"b7",  x"22",  x"82",  x"b7",  x"13", -- 25E0
         x"cd",  x"03",  x"f0",  x"18",  x"38",  x"d1",  x"2a",  x"97", -- 25E8
         x"b7",  x"22",  x"84",  x"b7",  x"13",  x"cd",  x"03",  x"f0", -- 25F0
         x"18",  x"38",  x"c4",  x"3a",  x"96",  x"b7",  x"b7",  x"67", -- 25F8
         x"6f",  x"28",  x"09",  x"2a",  x"97",  x"b7",  x"ed",  x"5b", -- 2600
         x"82",  x"b7",  x"ed",  x"52",  x"22",  x"f5",  x"b7",  x"3e", -- 2608
         x"0a",  x"cd",  x"13",  x"cb",  x"cd",  x"03",  x"f0",  x"23", -- 2610
         x"02",  x"4d",  x"61",  x"72",  x"6b",  x"65",  x"6e",  x"62", -- 2618
         x"65",  x"72",  x"65",  x"69",  x"63",  x"68",  x"3a",  x"20", -- 2620
         x"00",  x"2a",  x"82",  x"b7",  x"ed",  x"5b",  x"84",  x"b7", -- 2628
         x"cd",  x"03",  x"f0",  x"1b",  x"01",  x"17",  x"0f",  x"cd", -- 2630
         x"3d",  x"cf",  x"d8",  x"cd",  x"03",  x"f0",  x"18",  x"38", -- 2638
         x"d3",  x"2a",  x"97",  x"b7",  x"22",  x"86",  x"b7",  x"13", -- 2640
         x"cd",  x"03",  x"f0",  x"18",  x"38",  x"c6",  x"2a",  x"97", -- 2648
         x"b7",  x"22",  x"88",  x"b7",  x"3e",  x"0a",  x"cd",  x"13", -- 2650
         x"cb",  x"cd",  x"e9",  x"cf",  x"21",  x"00",  x"02",  x"24", -- 2658
         x"7c",  x"fe",  x"c0",  x"28",  x"08",  x"7e",  x"2f",  x"77", -- 2660
         x"be",  x"2f",  x"77",  x"28",  x"f2",  x"22",  x"80",  x"a8", -- 2668
         x"cd",  x"e0",  x"cf",  x"2a",  x"80",  x"a8",  x"cd",  x"03", -- 2670
         x"f0",  x"23",  x"02",  x"4d",  x"61",  x"72",  x"6b",  x"65", -- 2678
         x"6e",  x"74",  x"61",  x"62",  x"65",  x"6c",  x"6c",  x"65", -- 2680
         x"3a",  x"20",  x"00",  x"cd",  x"03",  x"f0",  x"1a",  x"01", -- 2688
         x"12",  x"0f",  x"cd",  x"3d",  x"cf",  x"d8",  x"cd",  x"03", -- 2690
         x"f0",  x"18",  x"38",  x"d7",  x"2a",  x"97",  x"b7",  x"22", -- 2698
         x"80",  x"a8",  x"cd",  x"03",  x"f0",  x"23",  x"0a",  x"02", -- 26A0
         x"4d",  x"61",  x"72",  x"6b",  x"65",  x"6e",  x"73",  x"63", -- 26A8
         x"68",  x"61",  x"6c",  x"74",  x"65",  x"72",  x"3a",  x"00", -- 26B0
         x"21",  x"f2",  x"b7",  x"36",  x"00",  x"3e",  x"10",  x"32", -- 26B8
         x"a0",  x"b7",  x"cb",  x"66",  x"28",  x"0a",  x"cd",  x"03", -- 26C0
         x"f0",  x"23",  x"45",  x"49",  x"4e",  x"00",  x"18",  x"08", -- 26C8
         x"cd",  x"03",  x"f0",  x"23",  x"41",  x"55",  x"53",  x"00", -- 26D0
         x"cd",  x"03",  x"f0",  x"04",  x"fe",  x"03",  x"c8",  x"fe", -- 26D8
         x"0d",  x"28",  x"0a",  x"fe",  x"20",  x"20",  x"f1",  x"3e", -- 26E0
         x"10",  x"ae",  x"77",  x"18",  x"d0",  x"cd",  x"03",  x"f0", -- 26E8
         x"23",  x"0a",  x"02",  x"50",  x"72",  x"6f",  x"6c",  x"6f", -- 26F0
         x"67",  x"62",  x"79",  x"74",  x"65",  x"73",  x"3a",  x"0d", -- 26F8
         x"0a",  x"00",  x"3e",  x"02",  x"cd",  x"03",  x"f0",  x"00", -- 2700
         x"06",  x"04",  x"21",  x"86",  x"c3",  x"7e",  x"cd",  x"03", -- 2708
         x"f0",  x"1c",  x"3e",  x"20",  x"cd",  x"13",  x"cb",  x"23", -- 2710
         x"10",  x"f3",  x"01",  x"12",  x"00",  x"cd",  x"3d",  x"cf", -- 2718
         x"d8",  x"06",  x"06",  x"21",  x"f7",  x"b7",  x"e5",  x"cd", -- 2720
         x"03",  x"f0",  x"18",  x"e1",  x"38",  x"d4",  x"3a",  x"97", -- 2728
         x"b7",  x"77",  x"13",  x"23",  x"10",  x"f0",  x"cd",  x"03", -- 2730
         x"f0",  x"23",  x"0a",  x"02",  x"32",  x"2e",  x"54",  x"72", -- 2738
         x"65",  x"6e",  x"6e",  x"7a",  x"65",  x"69",  x"63",  x"68", -- 2740
         x"65",  x"6e",  x"3a",  x"00",  x"21",  x"f2",  x"b7",  x"3e", -- 2748
         x"10",  x"32",  x"a0",  x"b7",  x"cb",  x"76",  x"28",  x"0a", -- 2750
         x"cd",  x"03",  x"f0",  x"23",  x"53",  x"50",  x"43",  x"00", -- 2758
         x"18",  x"08",  x"cd",  x"03",  x"f0",  x"23",  x"54",  x"41", -- 2760
         x"42",  x"00",  x"cd",  x"03",  x"f0",  x"04",  x"fe",  x"03", -- 2768
         x"c8",  x"fe",  x"0d",  x"28",  x"0a",  x"fe",  x"20",  x"20", -- 2770
         x"f1",  x"3e",  x"40",  x"ae",  x"77",  x"18",  x"d0",  x"cd", -- 2778
         x"03",  x"f0",  x"23",  x"0a",  x"02",  x"44",  x"65",  x"76", -- 2780
         x"69",  x"63",  x"65",  x"3d",  x"00",  x"3e",  x"fe",  x"cd", -- 2788
         x"03",  x"f0",  x"49",  x"cd",  x"03",  x"f0",  x"23",  x"2c", -- 2790
         x"20",  x"50",  x"72",  x"69",  x"6e",  x"74",  x"2c",  x"20", -- 2798
         x"53",  x"63",  x"72",  x"65",  x"65",  x"6e",  x"2c",  x"20", -- 27A0
         x"41",  x"73",  x"73",  x"65",  x"6d",  x"62",  x"6c",  x"65", -- 27A8
         x"72",  x"3f",  x"20",  x"00",  x"cd",  x"03",  x"f0",  x"04", -- 27B0
         x"fe",  x"03",  x"c8",  x"e6",  x"df",  x"2e",  x"01",  x"fe", -- 27B8
         x"44",  x"28",  x"0f",  x"2c",  x"fe",  x"50",  x"28",  x"0a", -- 27C0
         x"2c",  x"fe",  x"53",  x"28",  x"05",  x"2c",  x"fe",  x"41", -- 27C8
         x"20",  x"e2",  x"cd",  x"03",  x"f0",  x"00",  x"cd",  x"03", -- 27D0
         x"f0",  x"23",  x"0a",  x"02",  x"00",  x"26",  x"00",  x"22", -- 27D8
         x"f3",  x"b7",  x"3e",  x"04",  x"bd",  x"20",  x"43",  x"cd", -- 27E0
         x"03",  x"f0",  x"23",  x"02",  x"54",  x"6f",  x"70",  x"20", -- 27E8
         x"6f",  x"66",  x"20",  x"52",  x"41",  x"4d",  x"3a",  x"20", -- 27F0
         x"30",  x"32",  x"30",  x"30",  x"00",  x"01",  x"0f",  x"0c", -- 27F8
         x"cd",  x"3d",  x"cf",  x"d8",  x"cd",  x"03",  x"f0",  x"18", -- 2800
         x"38",  x"dd",  x"2a",  x"97",  x"b7",  x"22",  x"42",  x"00", -- 2808
         x"cd",  x"e9",  x"cf",  x"36",  x"0d",  x"cd",  x"e0",  x"cf", -- 2810
         x"23",  x"22",  x"18",  x"00",  x"22",  x"1c",  x"00",  x"2a", -- 2818
         x"80",  x"a8",  x"22",  x"46",  x"00",  x"22",  x"44",  x"00", -- 2820
         x"18",  x"3c",  x"3e",  x"02",  x"bd",  x"20",  x"3e",  x"cd", -- 2828
         x"03",  x"f0",  x"23",  x"02",  x"52",  x"61",  x"6e",  x"64", -- 2830
         x"20",  x"5a",  x"65",  x"69",  x"6c",  x"65",  x"6e",  x"3a", -- 2838
         x"20",  x"00",  x"01",  x"11",  x"0d",  x"cd",  x"3d",  x"cf", -- 2840
         x"d8",  x"cd",  x"03",  x"f0",  x"18",  x"38",  x"e0",  x"3a", -- 2848
         x"97",  x"b7",  x"32",  x"92",  x"b7",  x"13",  x"cd",  x"03", -- 2850
         x"f0",  x"18",  x"38",  x"d3",  x"3a",  x"97",  x"b7",  x"32", -- 2858
         x"93",  x"b7",  x"af",  x"32",  x"94",  x"b7",  x"cd",  x"03", -- 2860
         x"f0",  x"23",  x"0a",  x"02",  x"00",  x"cd",  x"03",  x"f0", -- 2868
         x"23",  x"0a",  x"02",  x"4f",  x"6b",  x"20",  x"3f",  x"20", -- 2870
         x"28",  x"4a",  x"29",  x"2f",  x"4e",  x"0a",  x"02",  x"00", -- 2878
         x"cd",  x"03",  x"f0",  x"04",  x"fe",  x"03",  x"c8",  x"e6", -- 2880
         x"df",  x"fe",  x"4e",  x"c8",  x"2a",  x"80",  x"a8",  x"2b", -- 2888
         x"22",  x"84",  x"a8",  x"cd",  x"03",  x"f0",  x"23",  x"0a", -- 2890
         x"02",  x"50",  x"41",  x"53",  x"53",  x"20",  x"31",  x"00", -- 2898
         x"cd",  x"bc",  x"cc",  x"3a",  x"f3",  x"b7",  x"fe",  x"04", -- 28A0
         x"20",  x"07",  x"2a",  x"82",  x"a8",  x"2b",  x"22",  x"1e", -- 28A8
         x"00",  x"cd",  x"03",  x"f0",  x"23",  x"08",  x"32",  x"0a", -- 28B0
         x"02",  x"00",  x"3a",  x"f3",  x"b7",  x"3d",  x"20",  x"2c", -- 28B8
         x"21",  x"e8",  x"c8",  x"cd",  x"ea",  x"ca",  x"d8",  x"21", -- 28C0
         x"00",  x"b7",  x"cd",  x"21",  x"f0",  x"02",  x"d8",  x"3e", -- 28C8
         x"02",  x"cd",  x"03",  x"f0",  x"00",  x"dd",  x"7e",  x"02", -- 28D0
         x"cd",  x"03",  x"f0",  x"1c",  x"3e",  x"3e",  x"cd",  x"03", -- 28D8
         x"f0",  x"00",  x"af",  x"32",  x"da",  x"b7",  x"18",  x"04", -- 28E0
         x"41",  x"53",  x"4d",  x"00",  x"af",  x"32",  x"91",  x"b7", -- 28E8
         x"21",  x"f2",  x"b7",  x"cb",  x"ae",  x"cd",  x"4f",  x"cb", -- 28F0
         x"cd",  x"4b",  x"cb",  x"3e",  x"4f",  x"cd",  x"56",  x"cb", -- 28F8
         x"3e",  x"52",  x"cd",  x"56",  x"cb",  x"3e",  x"47",  x"cd", -- 2900
         x"56",  x"cb",  x"cd",  x"42",  x"cb",  x"3e",  x"30",  x"cd", -- 2908
         x"56",  x"cb",  x"2a",  x"82",  x"b7",  x"cd",  x"7e",  x"c3", -- 2910
         x"cd",  x"24",  x"cb",  x"3e",  x"48",  x"cd",  x"56",  x"cb", -- 2918
         x"cd",  x"4f",  x"cb",  x"3e",  x"3b",  x"cd",  x"56",  x"cb", -- 2920
         x"cd",  x"03",  x"f0",  x"2a",  x"38",  x"4c",  x"21",  x"88", -- 2928
         x"a8",  x"22",  x"86",  x"a8",  x"11",  x"89",  x"a8",  x"01", -- 2930
         x"30",  x"00",  x"36",  x"00",  x"ed",  x"b0",  x"2a",  x"82", -- 2938
         x"b7",  x"ed",  x"5b",  x"84",  x"b7",  x"b7",  x"ed",  x"52", -- 2940
         x"d2",  x"7b",  x"ca",  x"3a",  x"f3",  x"b7",  x"fe",  x"04", -- 2948
         x"c2",  x"e0",  x"c9",  x"2a",  x"1e",  x"00",  x"ed",  x"5b", -- 2950
         x"1c",  x"00",  x"b7",  x"ed",  x"52",  x"d2",  x"e0",  x"c9", -- 2958
         x"cd",  x"03",  x"f0",  x"23",  x"0d",  x"0a",  x"3c",  x"3c", -- 2960
         x"3c",  x"20",  x"4e",  x"6f",  x"20",  x"4d",  x"65",  x"6d", -- 2968
         x"6f",  x"72",  x"79",  x"20",  x"3e",  x"3e",  x"3e",  x"0d", -- 2970
         x"0a",  x"00",  x"3a",  x"f3",  x"b7",  x"fe",  x"04",  x"20", -- 2978
         x"42",  x"cd",  x"e9",  x"cf",  x"2a",  x"1c",  x"00",  x"ed", -- 2980
         x"4b",  x"18",  x"00",  x"a7",  x"ed",  x"42",  x"44",  x"4d", -- 2988
         x"2a",  x"46",  x"00",  x"2b",  x"22",  x"1a",  x"00",  x"36", -- 2990
         x"03",  x"2b",  x"36",  x"0a",  x"2b",  x"36",  x"0d",  x"2b", -- 2998
         x"eb",  x"2a",  x"1c",  x"00",  x"2b",  x"ed",  x"b8",  x"23", -- 29A0
         x"22",  x"1c",  x"00",  x"13",  x"ed",  x"53",  x"1e",  x"00", -- 29A8
         x"ed",  x"43",  x"20",  x"00",  x"ed",  x"43",  x"40",  x"00", -- 29B0
         x"21",  x"08",  x"28",  x"22",  x"10",  x"00",  x"cd",  x"e0", -- 29B8
         x"cf",  x"18",  x"15",  x"cd",  x"4f",  x"cb",  x"3e",  x"03", -- 29C0
         x"cd",  x"56",  x"cb",  x"3a",  x"f3",  x"b7",  x"3d",  x"20", -- 29C8
         x"07",  x"01",  x"00",  x"01",  x"cd",  x"21",  x"f0",  x"03", -- 29D0
         x"cd",  x"03",  x"f0",  x"23",  x"0a",  x"02",  x"00",  x"c9", -- 29D8
         x"ed",  x"5b",  x"82",  x"b7",  x"3a",  x"f4",  x"b7",  x"f5", -- 29E0
         x"d5",  x"cd",  x"9c",  x"c3",  x"ed",  x"53",  x"82",  x"b7", -- 29E8
         x"21",  x"f2",  x"b7",  x"cb",  x"ee",  x"e1",  x"e5",  x"cd", -- 29F0
         x"4f",  x"cb",  x"cd",  x"7e",  x"c3",  x"cd",  x"7a",  x"cd", -- 29F8
         x"e1",  x"f1",  x"fe",  x"05",  x"28",  x"16",  x"b7",  x"20", -- 2A00
         x"6d",  x"cd",  x"d9",  x"cd",  x"28",  x"0e",  x"38",  x"0c", -- 2A08
         x"3a",  x"f2",  x"b7",  x"cb",  x"67",  x"28",  x"5f",  x"cd", -- 2A10
         x"ad",  x"ce",  x"20",  x"5a",  x"21",  x"88",  x"a8",  x"7e", -- 2A18
         x"fe",  x"30",  x"38",  x"04",  x"fe",  x"3a",  x"38",  x"06", -- 2A20
         x"cd",  x"56",  x"cb",  x"23",  x"18",  x"f1",  x"06",  x"05", -- 2A28
         x"e5",  x"7e",  x"b7",  x"28",  x"14",  x"fe",  x"48",  x"28", -- 2A30
         x"10",  x"fe",  x"2c",  x"28",  x"0c",  x"fe",  x"29",  x"28", -- 2A38
         x"08",  x"fe",  x"2d",  x"28",  x"04",  x"05",  x"23",  x"18", -- 2A40
         x"e8",  x"78",  x"a7",  x"20",  x"04",  x"e1",  x"23",  x"e5", -- 2A48
         x"3c",  x"47",  x"3e",  x"55",  x"cd",  x"56",  x"cb",  x"3e", -- 2A50
         x"30",  x"10",  x"f9",  x"e1",  x"7e",  x"23",  x"b7",  x"ca", -- 2A58
         x"28",  x"c9",  x"fe",  x"48",  x"28",  x"05",  x"cd",  x"56", -- 2A60
         x"cb",  x"18",  x"f1",  x"7e",  x"b7",  x"ca",  x"28",  x"c9", -- 2A68
         x"cd",  x"56",  x"cb",  x"23",  x"18",  x"f5",  x"21",  x"88", -- 2A70
         x"a8",  x"18",  x"f0",  x"ed",  x"5b",  x"80",  x"a8",  x"2a", -- 2A78
         x"82",  x"a8",  x"b7",  x"ed",  x"52",  x"d2",  x"7a",  x"c9", -- 2A80
         x"eb",  x"cd",  x"e9",  x"cf",  x"2b",  x"3e",  x"ff",  x"be", -- 2A88
         x"20",  x"0d",  x"2b",  x"be",  x"20",  x"08",  x"22",  x"80", -- 2A90
         x"a8",  x"cd",  x"e0",  x"cf",  x"18",  x"dd",  x"23",  x"56", -- 2A98
         x"2b",  x"5e",  x"cd",  x"e0",  x"cf",  x"22",  x"80",  x"a8", -- 2AA0
         x"21",  x"f2",  x"b7",  x"cb",  x"8e",  x"eb",  x"cd",  x"4f", -- 2AA8
         x"cb",  x"cd",  x"ac",  x"cd",  x"3e",  x"45",  x"cd",  x"56", -- 2AB0
         x"cb",  x"3e",  x"51",  x"cd",  x"56",  x"cb",  x"3e",  x"55", -- 2AB8
         x"cd",  x"56",  x"cb",  x"cd",  x"42",  x"cb",  x"3e",  x"30", -- 2AC0
         x"cd",  x"56",  x"cb",  x"cd",  x"24",  x"cb",  x"3e",  x"48", -- 2AC8
         x"cd",  x"56",  x"cb",  x"3a",  x"f3",  x"b7",  x"fe",  x"04", -- 2AD0
         x"20",  x"a1",  x"2a",  x"1e",  x"00",  x"ed",  x"5b",  x"1c", -- 2AD8
         x"00",  x"25",  x"b7",  x"ed",  x"52",  x"da",  x"60",  x"c9", -- 2AE0
         x"18",  x"91",  x"cd",  x"23",  x"cf",  x"d8",  x"eb",  x"11", -- 2AE8
         x"00",  x"b7",  x"01",  x"0b",  x"00",  x"ed",  x"b0",  x"cd", -- 2AF0
         x"57",  x"d2",  x"af",  x"12",  x"1c",  x"f8",  x"18",  x"fb", -- 2AF8
         x"3a",  x"f2",  x"b7",  x"cb",  x"77",  x"3e",  x"09",  x"28", -- 2B00
         x"02",  x"3e",  x"20",  x"f5",  x"3a",  x"f3",  x"b7",  x"a7", -- 2B08
         x"20",  x"06",  x"f1",  x"cd",  x"03",  x"f0",  x"24",  x"c9", -- 2B10
         x"f1",  x"e5",  x"2a",  x"86",  x"a8",  x"77",  x"23",  x"22", -- 2B18
         x"86",  x"a8",  x"e1",  x"c9",  x"f5",  x"7c",  x"cd",  x"2f", -- 2B20
         x"cb",  x"7d",  x"cd",  x"2f",  x"cb",  x"f1",  x"c9",  x"f5", -- 2B28
         x"1f",  x"1f",  x"1f",  x"1f",  x"cd",  x"38",  x"cb",  x"f1", -- 2B30
         x"e6",  x"0f",  x"c6",  x"90",  x"27",  x"ce",  x"40",  x"27", -- 2B38
         x"18",  x"14",  x"3a",  x"f2",  x"b7",  x"cb",  x"77",  x"3e", -- 2B40
         x"20",  x"20",  x"0b",  x"3e",  x"09",  x"18",  x"07",  x"3e", -- 2B48
         x"0d",  x"cd",  x"56",  x"cb",  x"3e",  x"0a",  x"c5",  x"d5", -- 2B50
         x"e5",  x"f5",  x"3a",  x"f3",  x"b7",  x"a7",  x"28",  x"3f", -- 2B58
         x"3d",  x"28",  x"43",  x"3d",  x"28",  x"69",  x"3d",  x"28", -- 2B60
         x"12",  x"2a",  x"1c",  x"00",  x"f1",  x"cd",  x"e9",  x"cf", -- 2B68
         x"77",  x"cd",  x"e0",  x"cf",  x"23",  x"22",  x"1c",  x"00", -- 2B70
         x"c3",  x"7f",  x"cc",  x"cd",  x"03",  x"f0",  x"0c",  x"fe", -- 2B78
         x"13",  x"20",  x"08",  x"cd",  x"03",  x"f0",  x"04",  x"fe", -- 2B80
         x"13",  x"28",  x"f8",  x"f1",  x"fe",  x"09",  x"20",  x"10", -- 2B88
         x"3e",  x"20",  x"cd",  x"13",  x"cb",  x"3a",  x"a0",  x"b7", -- 2B90
         x"e6",  x"07",  x"ca",  x"7f",  x"cc",  x"18",  x"f1",  x"f1", -- 2B98
         x"cd",  x"13",  x"cb",  x"c3",  x"7f",  x"cc",  x"f1",  x"57", -- 2BA0
         x"3a",  x"da",  x"b7",  x"26",  x"b7",  x"6f",  x"72",  x"3c", -- 2BA8
         x"e6",  x"7f",  x"32",  x"da",  x"b7",  x"c2",  x"7f",  x"cc", -- 2BB0
         x"01",  x"00",  x"01",  x"cd",  x"21",  x"f0",  x"00",  x"3e", -- 2BB8
         x"19",  x"cd",  x"03",  x"f0",  x"00",  x"dd",  x"7e",  x"02", -- 2BC0
         x"cd",  x"03",  x"f0",  x"1c",  x"c3",  x"7f",  x"cc",  x"f1", -- 2BC8
         x"fe",  x"03",  x"c4",  x"83",  x"cc",  x"fe",  x"0a",  x"c2", -- 2BD0
         x"7f",  x"cc",  x"3a",  x"93",  x"b7",  x"b7",  x"28",  x"31", -- 2BD8
         x"47",  x"3a",  x"94",  x"b7",  x"3c",  x"b8",  x"38",  x"29", -- 2BE0
         x"3e",  x"0c",  x"cd",  x"b0",  x"cc",  x"cd",  x"03",  x"f0", -- 2BE8
         x"23",  x"4e",  x"65",  x"78",  x"74",  x"20",  x"50",  x"61", -- 2BF0
         x"67",  x"65",  x"21",  x"00",  x"cd",  x"03",  x"f0",  x"04", -- 2BF8
         x"f5",  x"3e",  x"02",  x"cd",  x"03",  x"f0",  x"00",  x"f1", -- 2C00
         x"fe",  x"03",  x"20",  x"04",  x"cd",  x"03",  x"f0",  x"12", -- 2C08
         x"af",  x"32",  x"94",  x"b7",  x"3a",  x"92",  x"b7",  x"b7", -- 2C10
         x"28",  x"09",  x"3c",  x"47",  x"3e",  x"20",  x"cd",  x"b0", -- 2C18
         x"cc",  x"10",  x"f9",  x"af",  x"32",  x"95",  x"b7",  x"21", -- 2C20
         x"f2",  x"b7",  x"cb",  x"4e",  x"28",  x"4c",  x"ed",  x"5b", -- 2C28
         x"82",  x"b7",  x"e1",  x"e5",  x"cd",  x"24",  x"cb",  x"eb", -- 2C30
         x"ed",  x"52",  x"7d",  x"fe",  x"04",  x"38",  x"02",  x"3e", -- 2C38
         x"04",  x"47",  x"d5",  x"c5",  x"3e",  x"20",  x"cd",  x"b0", -- 2C40
         x"cc",  x"1a",  x"13",  x"cd",  x"2f",  x"cb",  x"10",  x"f4", -- 2C48
         x"c1",  x"c5",  x"3e",  x"05",  x"90",  x"47",  x"3e",  x"20", -- 2C50
         x"cd",  x"b0",  x"cc",  x"3e",  x"20",  x"cd",  x"b0",  x"cc", -- 2C58
         x"3e",  x"20",  x"cd",  x"b0",  x"cc",  x"10",  x"ef",  x"c1", -- 2C60
         x"d1",  x"1a",  x"13",  x"fe",  x"7f",  x"30",  x"04",  x"fe", -- 2C68
         x"20",  x"30",  x"02",  x"3e",  x"2e",  x"cd",  x"b0",  x"cc", -- 2C70
         x"10",  x"ef",  x"3e",  x"09",  x"cd",  x"83",  x"cc",  x"e1", -- 2C78
         x"d1",  x"c1",  x"c9",  x"f5",  x"fe",  x"09",  x"28",  x"05", -- 2C80
         x"cd",  x"b0",  x"cc",  x"18",  x"12",  x"3a",  x"95",  x"b7", -- 2C88
         x"06",  x"19",  x"b8",  x"38",  x"0c",  x"06",  x"21",  x"b8", -- 2C90
         x"38",  x"07",  x"06",  x"26",  x"b8",  x"38",  x"02",  x"f1", -- 2C98
         x"c9",  x"c5",  x"3e",  x"20",  x"cd",  x"b0",  x"cc",  x"3a", -- 2CA0
         x"95",  x"b7",  x"c1",  x"b8",  x"20",  x"f3",  x"18",  x"ef", -- 2CA8
         x"cd",  x"03",  x"f0",  x"02",  x"3a",  x"95",  x"b7",  x"3c", -- 2CB0
         x"32",  x"95",  x"b7",  x"c9",  x"2a",  x"80",  x"a8",  x"22", -- 2CB8
         x"82",  x"a8",  x"2a",  x"88",  x"b7",  x"ed",  x"5b",  x"86", -- 2CC0
         x"b7",  x"b7",  x"2b",  x"ed",  x"52",  x"d8",  x"21",  x"f2", -- 2CC8
         x"b7",  x"cb",  x"56",  x"28",  x"10",  x"cb",  x"96",  x"eb", -- 2CD0
         x"5e",  x"23",  x"56",  x"23",  x"22",  x"86",  x"b7",  x"19", -- 2CD8
         x"cd",  x"7e",  x"c3",  x"18",  x"42",  x"eb",  x"cd",  x"d9", -- 2CE0
         x"cd",  x"e5",  x"f5",  x"09",  x"22",  x"86",  x"b7",  x"21", -- 2CE8
         x"f2",  x"b7",  x"cb",  x"5e",  x"28",  x"04",  x"e1",  x"e1", -- 2CF0
         x"18",  x"c8",  x"f1",  x"e1",  x"28",  x"0e",  x"38",  x"18", -- 2CF8
         x"3a",  x"f2",  x"b7",  x"cb",  x"67",  x"28",  x"bb",  x"cd", -- 2D00
         x"ad",  x"ce",  x"20",  x"b6",  x"79",  x"fe",  x"04",  x"20", -- 2D08
         x"01",  x"23",  x"23",  x"5e",  x"23",  x"56",  x"18",  x"10", -- 2D10
         x"23",  x"7e",  x"23",  x"4f",  x"06",  x"00",  x"fe",  x"80", -- 2D18
         x"38",  x"01",  x"25",  x"09",  x"cd",  x"7e",  x"c3",  x"eb", -- 2D20
         x"2a",  x"82",  x"a8",  x"ed",  x"4b",  x"80",  x"a8",  x"e5", -- 2D28
         x"b7",  x"ed",  x"42",  x"e1",  x"30",  x"18",  x"cd",  x"e9", -- 2D30
         x"cf",  x"4e",  x"23",  x"46",  x"23",  x"cd",  x"e0",  x"cf", -- 2D38
         x"e5",  x"62",  x"6b",  x"b7",  x"ed",  x"42",  x"e1",  x"ca", -- 2D40
         x"c2",  x"cc",  x"38",  x"df",  x"2b",  x"2b",  x"ed",  x"4b", -- 2D48
         x"82",  x"a8",  x"c5",  x"d5",  x"cd",  x"e9",  x"cf",  x"50", -- 2D50
         x"59",  x"b7",  x"ed",  x"42",  x"28",  x"0a",  x"44",  x"4d", -- 2D58
         x"62",  x"6b",  x"1b",  x"1b",  x"ed",  x"b0",  x"13",  x"13", -- 2D60
         x"eb",  x"d1",  x"2b",  x"72",  x"2b",  x"73",  x"cd",  x"e0", -- 2D68
         x"cf",  x"e1",  x"2b",  x"2b",  x"22",  x"82",  x"a8",  x"c3", -- 2D70
         x"c2",  x"cc",  x"e5",  x"ed",  x"5b",  x"84",  x"a8",  x"2a", -- 2D78
         x"82",  x"a8",  x"2b",  x"b7",  x"ed",  x"52",  x"38",  x"07", -- 2D80
         x"e1",  x"cd",  x"e0",  x"cf",  x"c3",  x"4b",  x"cb",  x"cd", -- 2D88
         x"e9",  x"cf",  x"e1",  x"1a",  x"47",  x"1b",  x"1a",  x"4f", -- 2D90
         x"e5",  x"b7",  x"ed",  x"42",  x"e1",  x"28",  x"05",  x"38", -- 2D98
         x"e8",  x"1b",  x"18",  x"ef",  x"1b",  x"ed",  x"53",  x"84", -- 2DA0
         x"a8",  x"cd",  x"e0",  x"cf",  x"3e",  x"55",  x"cd",  x"56", -- 2DA8
         x"cb",  x"cd",  x"24",  x"cb",  x"cd",  x"4b",  x"cb",  x"ed", -- 2DB0
         x"5b",  x"84",  x"a8",  x"3e",  x"ff",  x"13",  x"cd",  x"e9", -- 2DB8
         x"cf",  x"12",  x"13",  x"12",  x"c3",  x"e0",  x"cf",  x"01", -- 2DC0
         x"02",  x"00",  x"3e",  x"1f",  x"23",  x"03",  x"be",  x"38", -- 2DC8
         x"fb",  x"21",  x"f2",  x"b7",  x"cb",  x"de",  x"c3",  x"8e", -- 2DD0
         x"ce",  x"e5",  x"d5",  x"3a",  x"f2",  x"b7",  x"e6",  x"f3", -- 2DD8
         x"32",  x"f2",  x"b7",  x"7e",  x"23",  x"be",  x"20",  x"10", -- 2DE0
         x"11",  x"f7",  x"b7",  x"06",  x"06",  x"4f",  x"1a",  x"b7", -- 2DE8
         x"28",  x"03",  x"b9",  x"28",  x"d2",  x"13",  x"10",  x"f6", -- 2DF0
         x"2b",  x"01",  x"04",  x"00",  x"7e",  x"fe",  x"ed",  x"28", -- 2DF8
         x"29",  x"cb",  x"af",  x"fe",  x"dd",  x"28",  x"09",  x"0d", -- 2E00
         x"7e",  x"fe",  x"cb",  x"20",  x"29",  x"0d",  x"18",  x"7e", -- 2E08
         x"23",  x"7e",  x"fe",  x"cb",  x"28",  x"78",  x"e6",  x"d8", -- 2E10
         x"fe",  x"30",  x"28",  x"0b",  x"7e",  x"e6",  x"c7",  x"fe", -- 2E18
         x"46",  x"28",  x"04",  x"fe",  x"86",  x"20",  x"0f",  x"0c", -- 2E20
         x"18",  x"0c",  x"23",  x"7e",  x"e6",  x"c7",  x"fe",  x"43", -- 2E28
         x"28",  x"5c",  x"0e",  x"02",  x"18",  x"58",  x"7e",  x"fe", -- 2E30
         x"cd",  x"28",  x"22",  x"fe",  x"c3",  x"28",  x"1b",  x"e6", -- 2E38
         x"e7",  x"fe",  x"22",  x"28",  x"49",  x"7e",  x"e6",  x"cf", -- 2E40
         x"fe",  x"01",  x"28",  x"42",  x"0d",  x"e6",  x"c7",  x"28", -- 2E48
         x"54",  x"fe",  x"c2",  x"28",  x"04",  x"fe",  x"c4",  x"20", -- 2E50
         x"39",  x"0c",  x"af",  x"18",  x"32",  x"23",  x"7e",  x"fe", -- 2E58
         x"21",  x"28",  x"04",  x"fe",  x"03",  x"20",  x"14",  x"23", -- 2E60
         x"7e",  x"fe",  x"f0",  x"20",  x"ed",  x"0c",  x"23",  x"7e", -- 2E68
         x"d6",  x"23",  x"20",  x"e6",  x"03",  x"23",  x"be",  x"20", -- 2E70
         x"fb",  x"18",  x"df",  x"fe",  x"0f",  x"20",  x"db",  x"23", -- 2E78
         x"7e",  x"fe",  x"f0",  x"20",  x"d5",  x"0e",  x"03",  x"21", -- 2E80
         x"f2",  x"b7",  x"cb",  x"d6",  x"18",  x"cc",  x"a7",  x"d1", -- 2E88
         x"e1",  x"c9",  x"fe",  x"06",  x"28",  x"f8",  x"fe",  x"c6", -- 2E90
         x"28",  x"f4",  x"7e",  x"e6",  x"f7",  x"fe",  x"d3",  x"28", -- 2E98
         x"ed",  x"0d",  x"79",  x"18",  x"e9",  x"7e",  x"fe",  x"09", -- 2EA0
         x"38",  x"f7",  x"37",  x"18",  x"e2",  x"e5",  x"c5",  x"d5", -- 2EA8
         x"cd",  x"d9",  x"cd",  x"79",  x"fe",  x"03",  x"30",  x"05", -- 2EB0
         x"d1",  x"c1",  x"e1",  x"a7",  x"c9",  x"7e",  x"fe",  x"dd", -- 2EB8
         x"28",  x"2f",  x"fe",  x"fd",  x"28",  x"2b",  x"fe",  x"ed", -- 2EC0
         x"28",  x"37",  x"fe",  x"01",  x"20",  x"05",  x"d1",  x"c1", -- 2EC8
         x"e1",  x"af",  x"c9",  x"fe",  x"11",  x"28",  x"f7",  x"fe", -- 2ED0
         x"21",  x"28",  x"f3",  x"fe",  x"31",  x"28",  x"ef",  x"fe", -- 2ED8
         x"22",  x"28",  x"eb",  x"fe",  x"2a",  x"28",  x"e7",  x"fe", -- 2EE0
         x"32",  x"28",  x"e3",  x"fe",  x"3a",  x"28",  x"df",  x"18", -- 2EE8
         x"c7",  x"23",  x"7e",  x"fe",  x"21",  x"28",  x"d7",  x"fe", -- 2EF0
         x"22",  x"28",  x"d3",  x"fe",  x"2a",  x"28",  x"cf",  x"18", -- 2EF8
         x"b7",  x"23",  x"7e",  x"fe",  x"43",  x"28",  x"c7",  x"fe", -- 2F00
         x"53",  x"28",  x"c3",  x"fe",  x"73",  x"28",  x"bf",  x"fe", -- 2F08
         x"4b",  x"28",  x"bb",  x"fe",  x"5b",  x"28",  x"b7",  x"fe", -- 2F10
         x"7b",  x"28",  x"b3",  x"18",  x"9b",  x"f5",  x"cd",  x"57", -- 2F18
         x"d2",  x"f1",  x"c9",  x"cd",  x"03",  x"f0",  x"23",  x"4e", -- 2F20
         x"61",  x"6d",  x"65",  x"20",  x"3a",  x"20",  x"20",  x"20", -- 2F28
         x"20",  x"20",  x"20",  x"20",  x"20",  x"00",  x"cd",  x"03", -- 2F30
         x"f0",  x"45",  x"01",  x"10",  x"06",  x"78",  x"32",  x"a0", -- 2F38
         x"b7",  x"cd",  x"03",  x"f0",  x"16",  x"fe",  x"03",  x"37", -- 2F40
         x"28",  x"d3",  x"fe",  x"0d",  x"28",  x"27",  x"fe",  x"20", -- 2F48
         x"30",  x"10",  x"fe",  x"09",  x"28",  x"0c",  x"fe",  x"08", -- 2F50
         x"28",  x"08",  x"fe",  x"1f",  x"28",  x"04",  x"fe",  x"0f", -- 2F58
         x"20",  x"df",  x"cd",  x"13",  x"cb",  x"3a",  x"a0",  x"b7", -- 2F60
         x"b8",  x"30",  x"01",  x"78",  x"b9",  x"38",  x"01",  x"79", -- 2F68
         x"32",  x"a0",  x"b7",  x"18",  x"cc",  x"ed",  x"5b",  x"a0", -- 2F70
         x"b7",  x"58",  x"cd",  x"03",  x"f0",  x"32",  x"eb",  x"c9", -- 2F78
         x"dd",  x"36",  x"02",  x"00",  x"21",  x"00",  x"b7",  x"1e", -- 2F80
         x"0b",  x"01",  x"f3",  x"83",  x"ed",  x"a3",  x"04",  x"04", -- 2F88
         x"1d",  x"20",  x"f9",  x"16",  x"0b",  x"dd",  x"34",  x"02", -- 2F90
         x"21",  x"00",  x"b7",  x"01",  x"f2",  x"81",  x"1e",  x"80", -- 2F98
         x"ed",  x"a3",  x"04",  x"04",  x"1d",  x"20",  x"f9",  x"7a", -- 2FA0
         x"01",  x"f3",  x"80",  x"ed",  x"79",  x"c5",  x"3e",  x"01", -- 2FA8
         x"cd",  x"03",  x"f0",  x"14",  x"c1",  x"ed",  x"78",  x"cb", -- 2FB0
         x"47",  x"20",  x"f2",  x"a7",  x"cb",  x"7f",  x"c8",  x"04", -- 2FB8
         x"ed",  x"78",  x"cd",  x"03",  x"f0",  x"1c",  x"cd",  x"03", -- 2FC0
         x"f0",  x"19",  x"37",  x"c9",  x"16",  x"03",  x"18",  x"c5", -- 2FC8
         x"cd",  x"cc",  x"cf",  x"d8",  x"16",  x"43",  x"dd",  x"36", -- 2FD0
         x"05",  x"00",  x"dd",  x"36",  x"06",  x"b7",  x"18",  x"c7", -- 2FD8
         x"f5",  x"db",  x"88",  x"f6",  x"24",  x"d3",  x"88",  x"f1", -- 2FE0
         x"c9",  x"f5",  x"db",  x"88",  x"e6",  x"db",  x"d3",  x"88", -- 2FE8
         x"f1",  x"c9",  x"e3",  x"2b",  x"e3",  x"e5",  x"f5",  x"2a", -- 2FF0
         x"a6",  x"00",  x"3a",  x"a8",  x"00",  x"77",  x"f1",  x"21", -- 2FF8
         x"6e",  x"d5",  x"18",  x"04",  x"e5",  x"21",  x"7f",  x"d5", -- 3000
         x"e3",  x"f5",  x"e5",  x"d5",  x"c5",  x"11",  x"28",  x"00", -- 3008
         x"21",  x"2c",  x"00",  x"01",  x"04",  x"00",  x"ed",  x"b0", -- 3010
         x"21",  x"0a",  x"00",  x"39",  x"7e",  x"23",  x"66",  x"6f", -- 3018
         x"0e",  x"0a",  x"ed",  x"b0",  x"c1",  x"d1",  x"e1",  x"db", -- 3020
         x"88",  x"f5",  x"3e",  x"8f",  x"d3",  x"88",  x"f1",  x"32", -- 3028
         x"8f",  x"00",  x"dd",  x"7e",  x"04",  x"32",  x"88",  x"00", -- 3030
         x"3e",  x"43",  x"dd",  x"77",  x"04",  x"d3",  x"86",  x"f1", -- 3038
         x"c9",  x"3e",  x"43",  x"dd",  x"77",  x"04",  x"d3",  x"86", -- 3040
         x"3e",  x"8f",  x"d3",  x"88",  x"3a",  x"a9",  x"00",  x"a7", -- 3048
         x"28",  x"0c",  x"3e",  x"87",  x"f3",  x"d3",  x"8c",  x"3e", -- 3050
         x"02",  x"d3",  x"8c",  x"fb",  x"00",  x"00",  x"f1",  x"c9", -- 3058
         x"fd",  x"fd",  x"57",  x"4f",  x"52",  x"4b",  x"52",  x"41", -- 3060
         x"4d",  x"01",  x"3d",  x"7d",  x"28",  x"02",  x"3e",  x"01", -- 3068
         x"cd",  x"03",  x"f0",  x"31",  x"cd",  x"49",  x"d7",  x"dd", -- 3070
         x"36",  x"09",  x"fd",  x"18",  x"3a",  x"7f",  x"7f",  x"54", -- 3078
         x"45",  x"4d",  x"4f",  x"01",  x"21",  x"10",  x"00",  x"af", -- 3080
         x"06",  x"18",  x"77",  x"23",  x"10",  x"fc",  x"21",  x"a6", -- 3088
         x"00",  x"06",  x"03",  x"77",  x"23",  x"10",  x"fc",  x"11", -- 3090
         x"e8",  x"aa",  x"21",  x"b0",  x"d1",  x"01",  x"0a",  x"00", -- 3098
         x"ed",  x"b0",  x"21",  x"a6",  x"b7",  x"ed",  x"a0",  x"ed", -- 30A0
         x"a0",  x"21",  x"86",  x"c3",  x"11",  x"f7",  x"b7",  x"01", -- 30A8
         x"06",  x"00",  x"ed",  x"b0",  x"cd",  x"46",  x"d7",  x"ed", -- 30B0
         x"57",  x"67",  x"2e",  x"60",  x"22",  x"24",  x"00",  x"2e", -- 30B8
         x"c4",  x"22",  x"ae",  x"b7",  x"f9",  x"dd",  x"22",  x"18", -- 30C0
         x"00",  x"af",  x"32",  x"81",  x"b7",  x"18",  x"22",  x"7f", -- 30C8
         x"7f",  x"52",  x"45",  x"54",  x"45",  x"4d",  x"4f",  x"01", -- 30D0
         x"ed",  x"57",  x"67",  x"2e",  x"c4",  x"22",  x"ae",  x"b7", -- 30D8
         x"f9",  x"cd",  x"46",  x"d7",  x"cd",  x"03",  x"f0",  x"12", -- 30E0
         x"fd",  x"fd",  x"4d",  x"45",  x"4e",  x"55",  x"01",  x"e1", -- 30E8
         x"e1",  x"cd",  x"03",  x"f0",  x"23",  x"1b",  x"32",  x"0c", -- 30F0
         x"0a",  x"3e",  x"20",  x"4b",  x"43",  x"2d",  x"44",  x"45", -- 30F8
         x"42",  x"55",  x"47",  x"47",  x"45",  x"52",  x"20",  x"32", -- 3100
         x"2e",  x"32",  x"20",  x"3c",  x"0d",  x"0a",  x"00",  x"cd", -- 3108
         x"03",  x"f0",  x"46",  x"2a",  x"a0",  x"b7",  x"22",  x"ed", -- 3110
         x"aa",  x"21",  x"f4",  x"aa",  x"ed",  x"4b",  x"36",  x"00", -- 3118
         x"79",  x"18",  x"2b",  x"11",  x"f4",  x"aa",  x"21",  x"9b", -- 3120
         x"b7",  x"01",  x"09",  x"00",  x"ed",  x"b0",  x"dd",  x"7e", -- 3128
         x"01",  x"e6",  x"0f",  x"12",  x"13",  x"23",  x"23",  x"ed", -- 3130
         x"a0",  x"ed",  x"a0",  x"21",  x"e8",  x"aa",  x"dd",  x"7e", -- 3138
         x"09",  x"32",  x"37",  x"00",  x"3a",  x"ec",  x"b7",  x"32", -- 3140
         x"36",  x"00",  x"3e",  x"2b",  x"06",  x"fd",  x"32",  x"ec", -- 3148
         x"b7",  x"dd",  x"70",  x"09",  x"11",  x"9b",  x"b7",  x"01", -- 3150
         x"09",  x"00",  x"ed",  x"b0",  x"3e",  x"1b",  x"cd",  x"13", -- 3158
         x"cb",  x"dd",  x"7e",  x"01",  x"e6",  x"f0",  x"b6",  x"dd", -- 3160
         x"77",  x"01",  x"d3",  x"84",  x"23",  x"13",  x"13",  x"ed", -- 3168
         x"a0",  x"ed",  x"a0",  x"e6",  x"01",  x"c6",  x"31",  x"c3", -- 3170
         x"13",  x"cb",  x"46",  x"20",  x"41",  x"20",  x"43",  x"20", -- 3178
         x"42",  x"20",  x"45",  x"20",  x"44",  x"20",  x"4c",  x"20", -- 3180
         x"48",  x"20",  x"53",  x"20",  x"5a",  x"20",  x"20",  x"20", -- 3188
         x"48",  x"59",  x"20",  x"20",  x"50",  x"20",  x"4e",  x"20", -- 3190
         x"43",  x"59",  x"41",  x"46",  x"42",  x"43",  x"44",  x"45", -- 3198
         x"48",  x"4c",  x"49",  x"59",  x"53",  x"50",  x"50",  x"43", -- 31A0
         x"53",  x"5a",  x"2e",  x"48",  x"2e",  x"50",  x"4e",  x"43", -- 31A8
         x"00",  x"00",  x"00",  x"28",  x"20",  x"00",  x"00",  x"00", -- 31B0
         x"39",  x"0d",  x"fd",  x"fd",  x"51",  x"55",  x"49",  x"54", -- 31B8
         x"01",  x"cd",  x"13",  x"d1",  x"ed",  x"57",  x"67",  x"2e", -- 31C0
         x"c4",  x"22",  x"ae",  x"b7",  x"f9",  x"cd",  x"03",  x"f0", -- 31C8
         x"12",  x"fd",  x"fd",  x"44",  x"49",  x"53",  x"41",  x"53", -- 31D0
         x"53",  x"01",  x"c3",  x"8d",  x"c4",  x"fd",  x"fd",  x"43", -- 31D8
         x"52",  x"43",  x"01",  x"fe",  x"02",  x"30",  x"19",  x"cd", -- 31E0
         x"03",  x"f0",  x"23",  x"0b",  x"09",  x"43",  x"52",  x"43", -- 31E8
         x"20",  x"41",  x"41",  x"44",  x"52",  x"20",  x"45",  x"41", -- 31F0
         x"44",  x"52",  x"2b",  x"31",  x"0d",  x"0a",  x"00",  x"c9", -- 31F8
         x"cd",  x"03",  x"d4",  x"11",  x"00",  x"00",  x"d5",  x"11", -- 3200
         x"ff",  x"ff",  x"7e",  x"e3",  x"85",  x"6f",  x"30",  x"01", -- 3208
         x"24",  x"e3",  x"7e",  x"aa",  x"57",  x"0f",  x"0f",  x"0f", -- 3210
         x"0f",  x"e6",  x"0f",  x"aa",  x"57",  x"0f",  x"0f",  x"0f", -- 3218
         x"f5",  x"e6",  x"1f",  x"ab",  x"5f",  x"f1",  x"f5",  x"0f", -- 3220
         x"e6",  x"f0",  x"ab",  x"5f",  x"f1",  x"e6",  x"e0",  x"aa", -- 3228
         x"53",  x"5f",  x"ed",  x"a1",  x"ea",  x"0a",  x"d2",  x"e1", -- 3230
         x"cd",  x"03",  x"f0",  x"23",  x"53",  x"55",  x"4d",  x"4d", -- 3238
         x"45",  x"3d",  x"00",  x"cd",  x"03",  x"f0",  x"1a",  x"eb", -- 3240
         x"cd",  x"03",  x"f0",  x"23",  x"43",  x"52",  x"43",  x"31", -- 3248
         x"36",  x"3d",  x"00",  x"cd",  x"03",  x"f0",  x"1a",  x"cd", -- 3250
         x"03",  x"f0",  x"2c",  x"c9",  x"fd",  x"fd",  x"52",  x"45", -- 3258
         x"47",  x"1f",  x"1a",  x"e6",  x"df",  x"ca",  x"ee",  x"d2", -- 3260
         x"21",  x"7a",  x"d1",  x"01",  x"2e",  x"00",  x"1a",  x"ed", -- 3268
         x"a1",  x"28",  x"07",  x"ed",  x"a1",  x"e2",  x"98",  x"d2", -- 3270
         x"18",  x"f4",  x"13",  x"1a",  x"fe",  x"40",  x"0b",  x"38", -- 3278
         x"09",  x"03",  x"ed",  x"a1",  x"1b",  x"20",  x"ee",  x"13", -- 3280
         x"13",  x"1a",  x"fe",  x"27",  x"20",  x"03",  x"13",  x"cb", -- 3288
         x"c0",  x"13",  x"cd",  x"03",  x"f0",  x"18",  x"30",  x"05", -- 3290
         x"cd",  x"03",  x"f0",  x"19",  x"c9",  x"ed",  x"5b",  x"97", -- 3298
         x"b7",  x"21",  x"10",  x"00",  x"3e",  x"2c",  x"91",  x"cb", -- 32A0
         x"6f",  x"20",  x"28",  x"0f",  x"cb",  x"5f",  x"28",  x"18", -- 32A8
         x"cb",  x"40",  x"28",  x"02",  x"2e",  x"1c",  x"e6",  x"07", -- 32B0
         x"01",  x"f8",  x"fd",  x"81",  x"4f",  x"0a",  x"cb",  x"43", -- 32B8
         x"28",  x"02",  x"b6",  x"01",  x"2f",  x"a6",  x"77",  x"c9", -- 32C0
         x"cb",  x"40",  x"28",  x"02",  x"c6",  x"0c",  x"c6",  x"10", -- 32C8
         x"6f",  x"73",  x"c9",  x"cb",  x"af",  x"2e",  x"1a",  x"fe", -- 32D0
         x"08",  x"28",  x"0f",  x"2e",  x"24",  x"fe",  x"0a",  x"28", -- 32D8
         x"09",  x"2e",  x"2a",  x"fe",  x"0c",  x"28",  x"03",  x"cd", -- 32E0
         x"c8",  x"d2",  x"73",  x"23",  x"72",  x"c9",  x"2a",  x"24", -- 32E8
         x"00",  x"7e",  x"23",  x"66",  x"6f",  x"22",  x"26",  x"00", -- 32F0
         x"cd",  x"03",  x"f0",  x"23",  x"41",  x"20",  x"20",  x"2d", -- 32F8
         x"46",  x"4c",  x"41",  x"47",  x"53",  x"2d",  x"2d",  x"20", -- 3300
         x"42",  x"20",  x"43",  x"20",  x"20",  x"44",  x"20",  x"45", -- 3308
         x"20",  x"20",  x"48",  x"20",  x"4c",  x"20",  x"20",  x"4d", -- 3310
         x"20",  x"20",  x"49",  x"58",  x"20",  x"20",  x"20",  x"49", -- 3318
         x"59",  x"20",  x"20",  x"20",  x"00",  x"21",  x"10",  x"00", -- 3320
         x"cd",  x"58",  x"d3",  x"cd",  x"03",  x"f0",  x"23",  x"41", -- 3328
         x"27",  x"20",  x"2d",  x"46",  x"4c",  x"41",  x"47",  x"53", -- 3330
         x"27",  x"2d",  x"20",  x"42",  x"27",  x"43",  x"27",  x"20", -- 3338
         x"44",  x"27",  x"45",  x"27",  x"20",  x"48",  x"27",  x"4c", -- 3340
         x"27",  x"20",  x"4d",  x"27",  x"20",  x"53",  x"50",  x"20", -- 3348
         x"20",  x"20",  x"28",  x"53",  x"50",  x"29",  x"20",  x"00", -- 3350
         x"4e",  x"23",  x"7e",  x"23",  x"cd",  x"d1",  x"d3",  x"06", -- 3358
         x"09",  x"11",  x"a8",  x"d1",  x"3e",  x"20",  x"cb",  x"21", -- 3360
         x"30",  x"01",  x"1a",  x"13",  x"cd",  x"13",  x"cb",  x"10", -- 3368
         x"f3",  x"06",  x"03",  x"cd",  x"7c",  x"d3",  x"1a",  x"cd", -- 3370
         x"d1",  x"d3",  x"06",  x"02",  x"5e",  x"23",  x"56",  x"23", -- 3378
         x"eb",  x"cd",  x"03",  x"f0",  x"1a",  x"eb",  x"10",  x"f4", -- 3380
         x"c9",  x"fd",  x"fd",  x"53",  x"57",  x"49",  x"54",  x"43", -- 3388
         x"48",  x"01",  x"fe",  x"01",  x"38",  x"31",  x"f5",  x"28", -- 3390
         x"0b",  x"53",  x"2d",  x"ca",  x"98",  x"d2",  x"2d",  x"ca", -- 3398
         x"98",  x"d2",  x"2c",  x"2c",  x"cd",  x"03",  x"f0",  x"26", -- 33A0
         x"5f",  x"7d",  x"cd",  x"d1",  x"d3",  x"7c",  x"cd",  x"d1", -- 33A8
         x"d3",  x"7b",  x"cd",  x"03",  x"f0",  x"1c",  x"f1",  x"28", -- 33B0
         x"0b",  x"3e",  x"09",  x"cd",  x"03",  x"f0",  x"42",  x"7a", -- 33B8
         x"cd",  x"03",  x"f0",  x"1c",  x"c3",  x"57",  x"d2",  x"cd", -- 33C0
         x"03",  x"f0",  x"23",  x"1b",  x"36",  x"1b",  x"35",  x"00", -- 33C8
         x"c9",  x"cd",  x"03",  x"f0",  x"1c",  x"cd",  x"03",  x"f0", -- 33D0
         x"2b",  x"c9",  x"fd",  x"fd",  x"44",  x"49",  x"53",  x"50", -- 33D8
         x"4c",  x"41",  x"59",  x"03",  x"cd",  x"03",  x"f0",  x"3b", -- 33E0
         x"c9",  x"fd",  x"fd",  x"4d",  x"4f",  x"44",  x"49",  x"46", -- 33E8
         x"59",  x"03",  x"cd",  x"03",  x"f0",  x"2e",  x"c9",  x"fd", -- 33F0
         x"fd",  x"2e",  x"01",  x"2a",  x"24",  x"00",  x"3e",  x"02", -- 33F8
         x"5f",  x"18",  x"ef",  x"eb",  x"2b",  x"ed",  x"52",  x"38", -- 3400
         x"07",  x"23",  x"eb",  x"c5",  x"42",  x"4b",  x"d1",  x"c9", -- 3408
         x"e1",  x"cd",  x"03",  x"f0",  x"23",  x"49",  x"4e",  x"56", -- 3410
         x"41",  x"4c",  x"49",  x"44",  x"20",  x"52",  x"41",  x"4e", -- 3418
         x"47",  x"45",  x"07",  x"00",  x"c3",  x"57",  x"d2",  x"fd", -- 3420
         x"fd",  x"49",  x"4e",  x"01",  x"3d",  x"28",  x"11",  x"cd", -- 3428
         x"03",  x"f0",  x"23",  x"0b",  x"09",  x"49",  x"4e",  x"20", -- 3430
         x"50",  x"4f",  x"52",  x"54",  x"0d",  x"0a",  x"00",  x"c9", -- 3438
         x"44",  x"4d",  x"ed",  x"78",  x"cd",  x"03",  x"f0",  x"1c", -- 3440
         x"c3",  x"57",  x"d2",  x"fd",  x"fd",  x"4f",  x"55",  x"54", -- 3448
         x"01",  x"fe",  x"02",  x"30",  x"22",  x"cd",  x"03",  x"f0", -- 3450
         x"23",  x"0b",  x"09",  x"4f",  x"55",  x"54",  x"20",  x"50", -- 3458
         x"4f",  x"52",  x"54",  x"20",  x"42",  x"59",  x"54",  x"45", -- 3460
         x"20",  x"28",  x"42",  x"59",  x"54",  x"45",  x"20",  x"2e", -- 3468
         x"2e",  x"2e",  x"29",  x"0d",  x"0a",  x"00",  x"c9",  x"44", -- 3470
         x"4d",  x"21",  x"82",  x"b7",  x"3d",  x"c8",  x"23",  x"23", -- 3478
         x"56",  x"ed",  x"51",  x"18",  x"f7",  x"fd",  x"fd",  x"46", -- 3480
         x"49",  x"4c",  x"4c",  x"01",  x"d6",  x"02",  x"30",  x"25", -- 3488
         x"cd",  x"03",  x"f0",  x"23",  x"0b",  x"09",  x"46",  x"49", -- 3490
         x"4c",  x"4c",  x"20",  x"41",  x"41",  x"44",  x"52",  x"20", -- 3498
         x"45",  x"41",  x"44",  x"52",  x"2b",  x"31",  x"20",  x"28", -- 34A0
         x"42",  x"59",  x"54",  x"45",  x"20",  x"2e",  x"2e",  x"2e", -- 34A8
         x"29",  x"0d",  x"0a",  x"00",  x"c9",  x"cd",  x"03",  x"d4", -- 34B0
         x"eb",  x"21",  x"86",  x"b7",  x"b7",  x"20",  x"03",  x"3c", -- 34B8
         x"36",  x"00",  x"f5",  x"e5",  x"ed",  x"a0",  x"e2",  x"d1", -- 34C0
         x"d4",  x"23",  x"3d",  x"20",  x"f7",  x"e1",  x"f1",  x"18", -- 34C8
         x"f1",  x"e1",  x"f1",  x"c9",  x"fd",  x"fd",  x"45",  x"58", -- 34D0
         x"43",  x"48",  x"01",  x"fe",  x"03",  x"28",  x"1f",  x"cd", -- 34D8
         x"03",  x"f0",  x"23",  x"0b",  x"09",  x"45",  x"58",  x"43", -- 34E0
         x"48",  x"20",  x"41",  x"41",  x"44",  x"52",  x"20",  x"45", -- 34E8
         x"41",  x"44",  x"52",  x"2b",  x"31",  x"20",  x"41",  x"44", -- 34F0
         x"52",  x"32",  x"0d",  x"0a",  x"00",  x"c9",  x"cd",  x"03", -- 34F8
         x"d4",  x"1a",  x"ed",  x"a0",  x"2b",  x"77",  x"23",  x"ea", -- 3500
         x"01",  x"d5",  x"c9",  x"fd",  x"fd",  x"43",  x"4f",  x"50", -- 3508
         x"59",  x"01",  x"fe",  x"03",  x"28",  x"1f",  x"cd",  x"03", -- 3510
         x"f0",  x"23",  x"0b",  x"09",  x"43",  x"4f",  x"50",  x"59", -- 3518
         x"20",  x"41",  x"41",  x"44",  x"52",  x"20",  x"45",  x"41", -- 3520
         x"44",  x"52",  x"2b",  x"31",  x"20",  x"41",  x"44",  x"52", -- 3528
         x"32",  x"0d",  x"0a",  x"00",  x"c9",  x"cd",  x"03",  x"d4", -- 3530
         x"ed",  x"52",  x"19",  x"38",  x"03",  x"ed",  x"b0",  x"c9", -- 3538
         x"09",  x"eb",  x"09",  x"eb",  x"2b",  x"1b",  x"ed",  x"b8", -- 3540
         x"c9",  x"fd",  x"fd",  x"42",  x"52",  x"45",  x"41",  x"4b", -- 3548
         x"01",  x"11",  x"57",  x"d2",  x"d5",  x"b7",  x"28",  x"03", -- 3550
         x"22",  x"a6",  x"00",  x"cd",  x"03",  x"f0",  x"23",  x"42", -- 3558
         x"52",  x"45",  x"41",  x"4b",  x"3d",  x"00",  x"2a",  x"a6", -- 3560
         x"00",  x"cd",  x"03",  x"f0",  x"1a",  x"c9",  x"f5",  x"e5", -- 3568
         x"2a",  x"a6",  x"00",  x"3a",  x"a8",  x"00",  x"77",  x"3e", -- 3570
         x"03",  x"32",  x"a9",  x"00",  x"e1",  x"18",  x"08",  x"f5", -- 3578
         x"3e",  x"03",  x"d3",  x"8c",  x"cd",  x"de",  x"d5",  x"f1", -- 3580
         x"ed",  x"73",  x"24",  x"00",  x"f3",  x"31",  x"24",  x"00", -- 3588
         x"d9",  x"e5",  x"d5",  x"c5",  x"d9",  x"08",  x"f5",  x"08", -- 3590
         x"fd",  x"e5",  x"dd",  x"e5",  x"e5",  x"d5",  x"c5",  x"f5", -- 3598
         x"ed",  x"7b",  x"24",  x"00",  x"2a",  x"2a",  x"00",  x"22", -- 35A0
         x"28",  x"00",  x"e1",  x"ed",  x"73",  x"24",  x"00",  x"22", -- 35A8
         x"2a",  x"00",  x"eb",  x"e1",  x"22",  x"26",  x"00",  x"e5", -- 35B0
         x"fb",  x"cd",  x"03",  x"f0",  x"0e",  x"30",  x"04",  x"fe", -- 35B8
         x"13",  x"28",  x"10",  x"2a",  x"a6",  x"00",  x"ed",  x"52", -- 35C0
         x"28",  x"09",  x"3a",  x"a9",  x"00",  x"3d",  x"ca",  x"29", -- 35C8
         x"d6",  x"18",  x"05",  x"3e",  x"03",  x"32",  x"a9",  x"00", -- 35D0
         x"cd",  x"23",  x"d1",  x"c3",  x"6a",  x"d6",  x"fb",  x"ed", -- 35D8
         x"4d",  x"fd",  x"fd",  x"47",  x"4f",  x"01",  x"a7",  x"28", -- 35E0
         x"0b",  x"22",  x"2a",  x"00",  x"11",  x"2c",  x"00",  x"01", -- 35E8
         x"04",  x"00",  x"ed",  x"b0",  x"db",  x"89",  x"f6",  x"1f", -- 35F0
         x"d3",  x"89",  x"2a",  x"a6",  x"00",  x"7e",  x"32",  x"a8", -- 35F8
         x"00",  x"36",  x"ff",  x"7e",  x"3c",  x"28",  x"02",  x"3e", -- 3600
         x"01",  x"32",  x"a9",  x"00",  x"cd",  x"19",  x"d1",  x"2a", -- 3608
         x"22",  x"00",  x"ed",  x"5b",  x"20",  x"00",  x"ed",  x"4b", -- 3610
         x"1e",  x"00",  x"d9",  x"2a",  x"1c",  x"00",  x"e5",  x"f1", -- 3618
         x"08",  x"ed",  x"4b",  x"12",  x"00",  x"ed",  x"7b",  x"24", -- 3620
         x"00",  x"2a",  x"2a",  x"00",  x"e5",  x"2a",  x"10",  x"00", -- 3628
         x"e5",  x"fd",  x"2a",  x"1a",  x"00",  x"2a",  x"16",  x"00", -- 3630
         x"ed",  x"5b",  x"14",  x"00",  x"c3",  x"87",  x"00",  x"fd", -- 3638
         x"fd",  x"53",  x"54",  x"45",  x"50",  x"01",  x"ed",  x"5b", -- 3640
         x"a0",  x"b7",  x"ed",  x"53",  x"ed",  x"aa",  x"a7",  x"28", -- 3648
         x"03",  x"22",  x"2a",  x"00",  x"db",  x"89",  x"f6",  x"1f", -- 3650
         x"d3",  x"89",  x"3e",  x"03",  x"32",  x"a9",  x"00",  x"2a", -- 3658
         x"2a",  x"00",  x"11",  x"2c",  x"00",  x"01",  x"0a",  x"00", -- 3660
         x"ed",  x"b0",  x"ed",  x"7b",  x"ae",  x"b7",  x"cd",  x"03", -- 3668
         x"f0",  x"2d",  x"cd",  x"f8",  x"d2",  x"af",  x"32",  x"f2", -- 3670
         x"b7",  x"67",  x"6f",  x"22",  x"f3",  x"b7",  x"2a",  x"28", -- 3678
         x"00",  x"11",  x"28",  x"00",  x"ed",  x"52",  x"22",  x"f5", -- 3680
         x"b7",  x"cd",  x"8c",  x"c3",  x"3e",  x"1d",  x"32",  x"a0", -- 3688
         x"b7",  x"af",  x"32",  x"f4",  x"b7",  x"cd",  x"5b",  x"d5", -- 3690
         x"2a",  x"2a",  x"00",  x"11",  x"2c",  x"00",  x"a7",  x"ed", -- 3698
         x"52",  x"22",  x"f5",  x"b7",  x"06",  x"02",  x"3e",  x"11", -- 36A0
         x"32",  x"a3",  x"b7",  x"c5",  x"cd",  x"8c",  x"c3",  x"cd", -- 36A8
         x"57",  x"d2",  x"c1",  x"3e",  x"39",  x"10",  x"f1",  x"3a", -- 36B0
         x"a9",  x"00",  x"fe",  x"02",  x"ca",  x"0c",  x"d6",  x"cd", -- 36B8
         x"03",  x"f0",  x"23",  x"02",  x"20",  x"57",  x"45",  x"49", -- 36C0
         x"54",  x"45",  x"52",  x"20",  x"4d",  x"49",  x"54",  x"3a", -- 36C8
         x"20",  x"43",  x"52",  x"2c",  x"20",  x"4c",  x"46",  x"2c", -- 36D0
         x"20",  x"42",  x"52",  x"4b",  x"2c",  x"20",  x"47",  x"2c", -- 36D8
         x"20",  x"55",  x"2c",  x"20",  x"49",  x"2c",  x"20",  x"53", -- 36E0
         x"3f",  x"00",  x"cd",  x"03",  x"f0",  x"16",  x"e6",  x"df", -- 36E8
         x"fe",  x"55",  x"28",  x"3d",  x"fe",  x"03",  x"28",  x"1b", -- 36F0
         x"fe",  x"0d",  x"ca",  x"0c",  x"d6",  x"fe",  x"0a",  x"28", -- 36F8
         x"1b",  x"fe",  x"49",  x"28",  x"20",  x"fe",  x"47",  x"ca", -- 3700
         x"fa",  x"d5",  x"fe",  x"53",  x"20",  x"dc",  x"3e",  x"02", -- 3708
         x"c3",  x"09",  x"d6",  x"2a",  x"ed",  x"aa",  x"22",  x"a0", -- 3710
         x"b7",  x"c3",  x"e4",  x"d0",  x"cd",  x"60",  x"d7",  x"22", -- 3718
         x"a6",  x"00",  x"c3",  x"fa",  x"d5",  x"2a",  x"2a",  x"00", -- 3720
         x"22",  x"28",  x"00",  x"cd",  x"60",  x"d7",  x"c3",  x"51", -- 3728
         x"d6",  x"2a",  x"a0",  x"b7",  x"e5",  x"cd",  x"19",  x"d1", -- 3730
         x"cd",  x"03",  x"f0",  x"04",  x"cd",  x"23",  x"d1",  x"e1", -- 3738
         x"22",  x"a0",  x"b7",  x"c3",  x"ea",  x"d6",  x"cd",  x"23", -- 3740
         x"d1",  x"11",  x"38",  x"00",  x"21",  x"f2",  x"cf",  x"01", -- 3748
         x"6e",  x"00",  x"ed",  x"b0",  x"ed",  x"57",  x"67",  x"2e", -- 3750
         x"e8",  x"11",  x"4a",  x"00",  x"73",  x"23",  x"72",  x"c9", -- 3758
         x"21",  x"2c",  x"00",  x"cd",  x"d9",  x"cd",  x"3a",  x"f2", -- 3760
         x"b7",  x"cb",  x"57",  x"28",  x"02",  x"03",  x"03",  x"2a", -- 3768
         x"2a",  x"00",  x"09",  x"c9",  x"7f",  x"7f",  x"53",  x"54", -- 3770
         x"41",  x"43",  x"4b",  x"20",  x"01",  x"21",  x"02",  x"00", -- 3778
         x"cd",  x"92",  x"d7",  x"c3",  x"f3",  x"db",  x"fd",  x"fd", -- 3780
         x"53",  x"54",  x"41",  x"43",  x"4b",  x"20",  x"01",  x"21", -- 3788
         x"00",  x"00",  x"39",  x"cd",  x"03",  x"f0",  x"1a",  x"7e", -- 3790
         x"23",  x"66",  x"6f",  x"cd",  x"03",  x"f0",  x"1a",  x"c3", -- 3798
         x"57",  x"d2",  x"7f",  x"7f",  x"4a",  x"20",  x"03",  x"7d", -- 37A0
         x"1e",  x"27",  x"c3",  x"09",  x"f0",  x"a1",  x"a1",  x"4d", -- 37A8
         x"45",  x"4e",  x"55",  x"01",  x"c3",  x"e2",  x"d8",  x"a1", -- 37B0
         x"a1",  x"41",  x"44",  x"52",  x"03",  x"e5",  x"11",  x"82", -- 37B8
         x"db",  x"ed",  x"57",  x"47",  x"0e",  x"75",  x"3e",  x"01", -- 37C0
         x"cd",  x"e6",  x"da",  x"e1",  x"e5",  x"1a",  x"13",  x"cd", -- 37C8
         x"e0",  x"da",  x"e1",  x"22",  x"a0",  x"aa",  x"cd",  x"e7", -- 37D0
         x"d7",  x"cd",  x"c8",  x"da",  x"21",  x"28",  x"11",  x"22", -- 37D8
         x"9e",  x"b7",  x"21",  x"00",  x"0f",  x"18",  x"09",  x"21", -- 37E0
         x"28",  x"20",  x"22",  x"9e",  x"b7",  x"21",  x"00",  x"00", -- 37E8
         x"22",  x"9c",  x"b7",  x"c9",  x"a1",  x"a1",  x"57",  x"41", -- 37F0
         x"49",  x"54",  x"03",  x"25",  x"24",  x"20",  x"1e",  x"7d", -- 37F8
         x"e6",  x"0f",  x"fe",  x"0a",  x"30",  x"17",  x"67",  x"ad", -- 3800
         x"0f",  x"6f",  x"0f",  x"0f",  x"85",  x"84",  x"fe",  x"40", -- 3808
         x"30",  x"0b",  x"32",  x"a4",  x"aa",  x"cd",  x"e7",  x"d7", -- 3810
         x"cd",  x"9f",  x"da",  x"18",  x"bf",  x"cd",  x"03",  x"f0", -- 3818
         x"19",  x"c9",  x"a1",  x"a1",  x"53",  x"41",  x"56",  x"45", -- 3820
         x"01",  x"21",  x"79",  x"db",  x"cd",  x"ea",  x"ca",  x"d8", -- 3828
         x"1e",  x"10",  x"21",  x"07",  x"db",  x"0e",  x"17",  x"ed", -- 3830
         x"b0",  x"cd",  x"f9",  x"da",  x"2a",  x"a0",  x"aa",  x"22", -- 3838
         x"1b",  x"b7",  x"21",  x"00",  x"b7",  x"dd",  x"75",  x"05", -- 3840
         x"dd",  x"74",  x"06",  x"cd",  x"03",  x"f0",  x"08",  x"d8", -- 3848
         x"cd",  x"03",  x"f0",  x"23",  x"02",  x"30",  x"31",  x"00", -- 3850
         x"dd",  x"36",  x"05",  x"17",  x"01",  x"a0",  x"00",  x"cd", -- 3858
         x"03",  x"f0",  x"09",  x"cd",  x"57",  x"d2",  x"c9",  x"a1", -- 3860
         x"a1",  x"45",  x"44",  x"49",  x"54",  x"1f",  x"cd",  x"c6", -- 3868
         x"d9",  x"38",  x"aa",  x"18",  x"6e",  x"7f",  x"7f",  x"4a", -- 3870
         x"45",  x"44",  x"49",  x"54",  x"1f",  x"3a",  x"80",  x"b7", -- 3878
         x"32",  x"b1",  x"aa",  x"21",  x"a9",  x"d9",  x"e5",  x"2a", -- 3880
         x"f0",  x"b7",  x"22",  x"a0",  x"aa",  x"22",  x"a2",  x"aa", -- 3888
         x"cd",  x"05",  x"da",  x"cd",  x"c6",  x"d9",  x"38",  x"d9", -- 3890
         x"3d",  x"28",  x"05",  x"3e",  x"02",  x"32",  x"a4",  x"aa", -- 3898
         x"dd",  x"36",  x"09",  x"a1",  x"21",  x"ec",  x"b7",  x"7e", -- 38A0
         x"32",  x"b0",  x"aa",  x"36",  x"2e",  x"ed",  x"57",  x"67", -- 38A8
         x"2e",  x"e1",  x"7e",  x"fe",  x"e0",  x"38",  x"0a",  x"21", -- 38B0
         x"7d",  x"db",  x"01",  x"92",  x"05",  x"ed",  x"b3",  x"18", -- 38B8
         x"21",  x"cd",  x"03",  x"f0",  x"23",  x"02",  x"66",  x"72", -- 38C0
         x"65",  x"6d",  x"64",  x"65",  x"20",  x"4a",  x"6f",  x"79", -- 38C8
         x"73",  x"74",  x"69",  x"63",  x"6b",  x"2d",  x"49",  x"53", -- 38D0
         x"52",  x"21",  x"07",  x"0d",  x"0a",  x"00",  x"cd",  x"03", -- 38D8
         x"f0",  x"04",  x"af",  x"f5",  x"cd",  x"43",  x"da",  x"f1", -- 38E0
         x"3d",  x"3e",  x"00",  x"32",  x"81",  x"b7",  x"20",  x"6c", -- 38E8
         x"cd",  x"03",  x"f0",  x"23",  x"0d",  x"0a",  x"50",  x"6c", -- 38F0
         x"65",  x"61",  x"73",  x"65",  x"2c",  x"20",  x"73",  x"65", -- 38F8
         x"6c",  x"65",  x"63",  x"74",  x"20",  x"6f",  x"72",  x"20", -- 3900
         x"70",  x"72",  x"65",  x"73",  x"73",  x"20",  x"53",  x"54", -- 3908
         x"4f",  x"50",  x"00",  x"21",  x"1e",  x"db",  x"22",  x"f0", -- 3910
         x"b7",  x"0e",  x"03",  x"06",  x"00",  x"79",  x"32",  x"a1", -- 3918
         x"b7",  x"21",  x"a2",  x"aa",  x"09",  x"11",  x"00",  x"09", -- 3920
         x"cd",  x"18",  x"da",  x"e5",  x"11",  x"38",  x"00",  x"19", -- 3928
         x"30",  x"04",  x"cd",  x"03",  x"f0",  x"25",  x"cd",  x"03", -- 3930
         x"f0",  x"0e",  x"30",  x"f3",  x"e1",  x"57",  x"fe",  x"13", -- 3938
         x"28",  x"2e",  x"d6",  x"80",  x"fe",  x"0b",  x"38",  x"2c", -- 3940
         x"72",  x"0c",  x"cd",  x"15",  x"da",  x"79",  x"fe",  x"0e", -- 3948
         x"38",  x"cb",  x"3c",  x"32",  x"a1",  x"b7",  x"3e",  x"02", -- 3950
         x"cd",  x"03",  x"f0",  x"00",  x"21",  x"2a",  x"db",  x"22", -- 3958
         x"f0",  x"b7",  x"cd",  x"dc",  x"d7",  x"26",  x"00",  x"22", -- 3960
         x"a0",  x"b7",  x"e1",  x"e1",  x"cd",  x"03",  x"f0",  x"46", -- 3968
         x"0e",  x"0e",  x"18",  x"d6",  x"c6",  x"03",  x"4f",  x"dd", -- 3970
         x"7e",  x"0d",  x"3d",  x"ba",  x"38",  x"f9",  x"18",  x"ca", -- 3978
         x"a1",  x"a1",  x"51",  x"55",  x"49",  x"54",  x"01",  x"2a", -- 3980
         x"a2",  x"aa",  x"22",  x"f0",  x"b7",  x"cd",  x"e7",  x"d7", -- 3988
         x"3a",  x"b0",  x"aa",  x"32",  x"ec",  x"b7",  x"3e",  x"7f", -- 3990
         x"dd",  x"77",  x"09",  x"11",  x"74",  x"db",  x"21",  x"00", -- 3998
         x"c0",  x"45",  x"4d",  x"cd",  x"03",  x"f0",  x"1d",  x"23", -- 39A0
         x"e3",  x"ed",  x"5b",  x"b0",  x"aa",  x"3e",  x"02",  x"6f", -- 39A8
         x"1e",  x"26",  x"c3",  x"09",  x"f0",  x"a1",  x"a1",  x"4f", -- 39B0
         x"4b",  x"01",  x"2a",  x"a0",  x"aa",  x"22",  x"f0",  x"b7", -- 39B8
         x"eb",  x"cd",  x"f9",  x"da",  x"18",  x"c7",  x"01",  x"a5", -- 39C0
         x"aa",  x"1a",  x"a7",  x"28",  x"17",  x"fe",  x"20",  x"28", -- 39C8
         x"0e",  x"fe",  x"2c",  x"28",  x"23",  x"cd",  x"03",  x"f0", -- 39D0
         x"18",  x"d8",  x"3a",  x"97",  x"b7",  x"02",  x"03",  x"13", -- 39D8
         x"cb",  x"61",  x"28",  x"e5",  x"3e",  x"a6",  x"91",  x"38", -- 39E0
         x"07",  x"c0",  x"0b",  x"0a",  x"a7",  x"28",  x"0d",  x"03", -- 39E8
         x"af",  x"cb",  x"61",  x"c0",  x"02",  x"03",  x"18",  x"f9", -- 39F0
         x"13",  x"1a",  x"18",  x"e1",  x"21",  x"94",  x"aa",  x"22", -- 39F8
         x"a0",  x"aa",  x"21",  x"2a",  x"db",  x"d5",  x"11",  x"a4", -- 3A00
         x"aa",  x"01",  x"42",  x"db",  x"ed",  x"a0",  x"0a",  x"5f", -- 3A08
         x"a7",  x"20",  x"f9",  x"d1",  x"c9",  x"56",  x"1e",  x"42", -- 3A10
         x"c5",  x"e5",  x"21",  x"a0",  x"b7",  x"36",  x"0d",  x"01", -- 3A18
         x"3c",  x"03",  x"7a",  x"a7",  x"3e",  x"3e",  x"20",  x"02", -- 3A20
         x"1e",  x"2b",  x"cd",  x"09",  x"f0",  x"7a",  x"51",  x"4f", -- 3A28
         x"10",  x"f8",  x"7b",  x"fe",  x"42",  x"20",  x"07",  x"36", -- 3A30
         x"13",  x"79",  x"cd",  x"03",  x"f0",  x"1c",  x"36",  x"0e", -- 3A38
         x"e1",  x"c1",  x"c9",  x"cd",  x"e7",  x"d7",  x"cd",  x"03", -- 3A40
         x"f0",  x"23",  x"0c",  x"0a",  x"2a",  x"20",  x"4a",  x"4f", -- 3A48
         x"59",  x"53",  x"54",  x"49",  x"43",  x"4b",  x"2d",  x"45", -- 3A50
         x"44",  x"49",  x"54",  x"4f",  x"52",  x"20",  x"2a",  x"20", -- 3A58
         x"20",  x"20",  x"41",  x"64",  x"72",  x"3a",  x"20",  x"20", -- 3A60
         x"20",  x"20",  x"20",  x"20",  x"57",  x"61",  x"69",  x"74", -- 3A68
         x"3a",  x"0d",  x"0a",  x"0a",  x"00",  x"21",  x"a5",  x"aa", -- 3A70
         x"e5",  x"21",  x"43",  x"db",  x"06",  x"0b",  x"e5",  x"5e", -- 3A78
         x"cb",  x"3b",  x"16",  x"00",  x"19",  x"cd",  x"03",  x"f0", -- 3A80
         x"45",  x"e1",  x"7e",  x"23",  x"0f",  x"30",  x"ef",  x"e3", -- 3A88
         x"cd",  x"15",  x"da",  x"23",  x"e3",  x"cd",  x"03",  x"f0", -- 3A90
         x"2c",  x"10",  x"e3",  x"e1",  x"cd",  x"c8",  x"da",  x"2a", -- 3A98
         x"a0",  x"b7",  x"11",  x"25",  x"01",  x"ed",  x"53",  x"a0", -- 3AA0
         x"b7",  x"3a",  x"a4",  x"aa",  x"11",  x"0a",  x"2f",  x"14", -- 3AA8
         x"93",  x"30",  x"fc",  x"c6",  x"3a",  x"5f",  x"7a",  x"fe", -- 3AB0
         x"30",  x"20",  x"02",  x"3e",  x"20",  x"cd",  x"03",  x"f0", -- 3AB8
         x"00",  x"7b",  x"cd",  x"03",  x"f0",  x"00",  x"18",  x"12", -- 3AC0
         x"2a",  x"a0",  x"b7",  x"e5",  x"21",  x"1a",  x"01",  x"22", -- 3AC8
         x"a0",  x"b7",  x"2a",  x"a0",  x"aa",  x"cd",  x"03",  x"f0", -- 3AD0
         x"1a",  x"e1",  x"22",  x"a0",  x"b7",  x"c9",  x"3d",  x"c8", -- 3AD8
         x"eb",  x"4e",  x"23",  x"46",  x"23",  x"eb",  x"a7",  x"ed", -- 3AE0
         x"42",  x"eb",  x"4e",  x"23",  x"46",  x"23",  x"eb",  x"a7", -- 3AE8
         x"ed",  x"42",  x"30",  x"ea",  x"f1",  x"f1",  x"c3",  x"11", -- 3AF0
         x"d4",  x"01",  x"42",  x"db",  x"21",  x"a4",  x"aa",  x"ed", -- 3AF8
         x"a0",  x"0a",  x"6f",  x"a7",  x"20",  x"f9",  x"c9",  x"03", -- 3B00
         x"80",  x"01",  x"9c",  x"01",  x"80",  x"01",  x"21",  x"90", -- 3B08
         x"01",  x"11",  x"00",  x"00",  x"ed",  x"53",  x"f0",  x"b7", -- 3B10
         x"01",  x"0c",  x"00",  x"ed",  x"b0",  x"c9",  x"02",  x"83", -- 3B18
         x"82",  x"8a",  x"80",  x"86",  x"88",  x"85",  x"81",  x"87", -- 3B20
         x"89",  x"84",  x"02",  x"0b",  x"0a",  x"0d",  x"08",  x"00", -- 3B28
         x"00",  x"0d",  x"09",  x"00",  x"00",  x"20",  x"00",  x"a9", -- 3B30
         x"ae",  x"ac",  x"a6",  x"aa",  x"ad",  x"ab",  x"a5",  x"af", -- 3B38
         x"a7",  x"a8",  x"a4",  x"25",  x"2f",  x"3b",  x"45",  x"4c", -- 3B40
         x"55",  x"49",  x"16",  x"39",  x"1e",  x"35",  x"0e",  x"25", -- 3B48
         x"16",  x"21",  x"36",  x"30",  x"3d",  x"6c",  x"65",  x"66", -- 3B50
         x"74",  x"20",  x"00",  x"72",  x"69",  x"67",  x"68",  x"74", -- 3B58
         x"00",  x"2b",  x"64",  x"6f",  x"77",  x"6e",  x"00",  x"2b", -- 3B60
         x"75",  x"70",  x"00",  x"20",  x"2b",  x"66",  x"69",  x"72", -- 3B68
         x"65",  x"00",  x"32",  x"00",  x"4d",  x"45",  x"4e",  x"55", -- 3B70
         x"00",  x"4a",  x"4f",  x"59",  x"00",  x"e0",  x"cf",  x"ff", -- 3B78
         x"97",  x"c0",  x"8b",  x"00",  x"04",  x"75",  x"01",  x"8b", -- 3B80
         x"00",  x"f5",  x"7d",  x"3b",  x"28",  x"c5",  x"04",  x"0b", -- 3B88
         x"0d",  x"f5",  x"05",  x"0b",  x"40",  x"fd",  x"fd",  x"3f", -- 3B90
         x"1f",  x"cd",  x"59",  x"dd",  x"28",  x"15",  x"cd",  x"9b", -- 3B98
         x"dc",  x"1e",  x"19",  x"da",  x"09",  x"f0",  x"cd",  x"66", -- 3BA0
         x"dd",  x"2a",  x"3f",  x"05",  x"22",  x"ae",  x"b7",  x"cd", -- 3BA8
         x"90",  x"dc",  x"c9",  x"cd",  x"03",  x"f0",  x"23",  x"0b", -- 3BB0
         x"09",  x"3f",  x"20",  x"41",  x"75",  x"73",  x"64",  x"72", -- 3BB8
         x"75",  x"63",  x"6b",  x"0d",  x"0a",  x"00",  x"c9",  x"7f", -- 3BC0
         x"7f",  x"3f",  x"63",  x"1f",  x"cd",  x"99",  x"db",  x"18", -- 3BC8
         x"22",  x"7f",  x"7f",  x"3f",  x"69",  x"01",  x"2a",  x"99", -- 3BD0
         x"b7",  x"11",  x"08",  x"01",  x"a7",  x"ed",  x"52",  x"28", -- 3BD8
         x"12",  x"19",  x"ed",  x"53",  x"99",  x"b7",  x"e5",  x"21", -- 3BE0
         x"26",  x"df",  x"01",  x"28",  x"00",  x"ed",  x"b0",  x"e1", -- 3BE8
         x"22",  x"2c",  x"01",  x"ed",  x"5b",  x"7f",  x"b7",  x"c3", -- 3BF0
         x"ad",  x"d9",  x"08",  x"f5",  x"c5",  x"d5",  x"e5",  x"fd", -- 3BF8
         x"e5",  x"cd",  x"9b",  x"dc",  x"38",  x"42",  x"21",  x"50", -- 3C00
         x"dc",  x"22",  x"99",  x"b7",  x"dd",  x"7e",  x"01",  x"f5", -- 3C08
         x"cb",  x"8f",  x"cb",  x"df",  x"dd",  x"77",  x"01",  x"21", -- 3C10
         x"a2",  x"b7",  x"36",  x"12",  x"e6",  x"01",  x"c6",  x"31", -- 3C18
         x"cd",  x"03",  x"f0",  x"00",  x"21",  x"28",  x"03",  x"22", -- 3C20
         x"9e",  x"b7",  x"ed",  x"62",  x"22",  x"9c",  x"b7",  x"22", -- 3C28
         x"ea",  x"03",  x"cd",  x"27",  x"dd",  x"cd",  x"03",  x"f0", -- 3C30
         x"23",  x"12",  x"0c",  x"00",  x"cd",  x"48",  x"dd",  x"38", -- 3C38
         x"15",  x"28",  x"2b",  x"cd",  x"66",  x"dd",  x"18",  x"f4", -- 3C40
         x"3e",  x"07",  x"cd",  x"03",  x"f0",  x"00",  x"18",  x"38", -- 3C48
         x"31",  x"0b",  x"0a",  x"37",  x"18",  x"18",  x"11",  x"ea", -- 3C50
         x"03",  x"cd",  x"59",  x"dd",  x"01",  x"0d",  x"00",  x"21", -- 3C58
         x"8e",  x"b9",  x"70",  x"23",  x"22",  x"62",  x"05",  x"eb", -- 3C60
         x"ed",  x"b0",  x"dd",  x"cb",  x"08",  x"f6",  x"08",  x"21", -- 3C68
         x"11",  x"05",  x"11",  x"80",  x"b7",  x"01",  x"80",  x"00", -- 3C70
         x"ed",  x"b0",  x"eb",  x"37",  x"cd",  x"27",  x"dd",  x"f1", -- 3C78
         x"dd",  x"77",  x"01",  x"d3",  x"84",  x"cd",  x"90",  x"dc", -- 3C80
         x"fd",  x"e1",  x"e1",  x"d1",  x"c1",  x"f1",  x"08",  x"c9", -- 3C88
         x"fd",  x"e1",  x"d1",  x"7a",  x"53",  x"e1",  x"f9",  x"06", -- 3C90
         x"01",  x"18",  x"18",  x"dd",  x"7c",  x"87",  x"d8",  x"d6", -- 3C98
         x"06",  x"fe",  x"0e",  x"d8",  x"fd",  x"e1",  x"db",  x"88", -- 3CA0
         x"5f",  x"21",  x"00",  x"c0",  x"45",  x"39",  x"30",  x"02", -- 3CA8
         x"f6",  x"0a",  x"57",  x"d5",  x"3d",  x"f3",  x"d3",  x"88", -- 3CB0
         x"dd",  x"7e",  x"01",  x"f5",  x"e6",  x"f9",  x"f6",  x"02", -- 3CB8
         x"d3",  x"84",  x"cd",  x"00",  x"dd",  x"06",  x"06",  x"f1", -- 3CC0
         x"10",  x"fd",  x"d3",  x"84",  x"e1",  x"7c",  x"d3",  x"88", -- 3CC8
         x"fb",  x"cb",  x"22",  x"30",  x"19",  x"ed",  x"73",  x"0f", -- 3CD0
         x"0a",  x"31",  x"0f",  x"0a",  x"e5",  x"21",  x"bd",  x"de", -- 3CD8
         x"11",  x"a8",  x"04",  x"0e",  x"69",  x"ed",  x"b0",  x"21", -- 3CE0
         x"80",  x"b7",  x"0e",  x"80",  x"ed",  x"b0",  x"dd",  x"36", -- 3CE8
         x"0d",  x"00",  x"3e",  x"14",  x"cd",  x"03",  x"f0",  x"14", -- 3CF0
         x"cd",  x"03",  x"f0",  x"0e",  x"38",  x"f0",  x"fd",  x"e9", -- 3CF8
         x"21",  x"86",  x"c3",  x"e5",  x"21",  x"f1",  x"d3",  x"e5", -- 3D00
         x"21",  x"ed",  x"b0",  x"e5",  x"21",  x"d3",  x"86",  x"e5", -- 3D08
         x"ed",  x"62",  x"39",  x"dd",  x"7e",  x"04",  x"f5",  x"f6", -- 3D10
         x"80",  x"e5",  x"21",  x"00",  x"03",  x"11",  x"00",  x"b8", -- 3D18
         x"10",  x"01",  x"eb",  x"01",  x"11",  x"07",  x"c9",  x"2a", -- 3D20
         x"cb",  x"b7",  x"01",  x"78",  x"00",  x"cd",  x"40",  x"dd", -- 3D28
         x"21",  x"00",  x"a7",  x"0e",  x"18",  x"cd",  x"40",  x"dd", -- 3D30
         x"7e",  x"2f",  x"77",  x"68",  x"25",  x"f0",  x"18",  x"f3", -- 3D38
         x"30",  x"01",  x"eb",  x"ed",  x"b0",  x"d0",  x"eb",  x"c9", -- 3D40
         x"3e",  x"3f",  x"cd",  x"03",  x"f0",  x"24",  x"cd",  x"03", -- 3D48
         x"f0",  x"17",  x"d8",  x"1a",  x"fe",  x"3f",  x"20",  x"01", -- 3D50
         x"13",  x"1a",  x"a7",  x"c8",  x"fe",  x"21",  x"38",  x"f8", -- 3D58
         x"ed",  x"53",  x"92",  x"b7",  x"a7",  x"c9",  x"ed",  x"73", -- 3D60
         x"ae",  x"b7",  x"21",  x"fe",  x"04",  x"22",  x"b9",  x"b7", -- 3D68
         x"23",  x"22",  x"be",  x"b7",  x"21",  x"bd",  x"c0",  x"11", -- 3D70
         x"00",  x"03",  x"01",  x"62",  x"00",  x"cd",  x"b4",  x"04", -- 3D78
         x"21",  x"61",  x"03",  x"0e",  x"9f",  x"ed",  x"b0",  x"21", -- 3D80
         x"a7",  x"04",  x"22",  x"b0",  x"03",  x"2e",  x"7f",  x"22", -- 3D88
         x"56",  x"03",  x"cd",  x"a8",  x"04",  x"3d",  x"32",  x"fc", -- 3D90
         x"03",  x"32",  x"58",  x"03",  x"2a",  x"92",  x"b7",  x"11", -- 3D98
         x"62",  x"03",  x"d5",  x"cd",  x"23",  x"de",  x"e1",  x"cd", -- 3DA0
         x"bb",  x"04",  x"cd",  x"e9",  x"dd",  x"3a",  x"ae",  x"03", -- 3DA8
         x"a7",  x"20",  x"21",  x"cd",  x"cb",  x"04",  x"eb",  x"d5", -- 3DB0
         x"cd",  x"92",  x"de",  x"d1",  x"c6",  x"30",  x"20",  x"10", -- 3DB8
         x"cd",  x"03",  x"f0",  x"2b",  x"cd",  x"03",  x"f0",  x"1a", -- 3DC0
         x"cd",  x"03",  x"f0",  x"23",  x"08",  x"48",  x"20",  x"00", -- 3DC8
         x"eb",  x"cd",  x"d3",  x"04",  x"cd",  x"db",  x"04",  x"ed", -- 3DD0
         x"7b",  x"ae",  x"b7",  x"3a",  x"a0",  x"b7",  x"a7",  x"c8", -- 3DD8
         x"cd",  x"03",  x"f0",  x"23",  x"20",  x"0d",  x"0a",  x"00", -- 3DE0
         x"c9",  x"e5",  x"2a",  x"4a",  x"05",  x"22",  x"b9",  x"b7", -- 3DE8
         x"2a",  x"4f",  x"05",  x"22",  x"be",  x"b7",  x"e1",  x"c9", -- 3DF0
         x"fe",  x"41",  x"38",  x"5e",  x"04",  x"10",  x"5b",  x"e5", -- 3DF8
         x"d5",  x"eb",  x"cd",  x"03",  x"f0",  x"18",  x"eb",  x"d1", -- 3E00
         x"7e",  x"e6",  x"df",  x"d6",  x"48",  x"20",  x"50",  x"23", -- 3E08
         x"e3",  x"d5",  x"ed",  x"5b",  x"97",  x"b7",  x"06",  x"98", -- 3E10
         x"cd",  x"c3",  x"04",  x"d1",  x"01",  x"01",  x"00",  x"cd", -- 3E18
         x"26",  x"de",  x"e1",  x"01",  x"00",  x"00",  x"7b",  x"fe", -- 3E20
         x"ab",  x"d0",  x"7e",  x"a7",  x"c8",  x"fe",  x"22",  x"28", -- 3E28
         x"28",  x"cb",  x"41",  x"20",  x"25",  x"fe",  x"3a",  x"30", -- 3E30
         x"08",  x"fe",  x"30",  x"30",  x"bf",  x"fe",  x"20",  x"28", -- 3E38
         x"15",  x"d5",  x"c5",  x"11",  x"20",  x"c1",  x"06",  x"80", -- 3E40
         x"cd",  x"6c",  x"de",  x"ed",  x"5b",  x"0c",  x"e0",  x"dc", -- 3E48
         x"6c",  x"de",  x"c1",  x"d1",  x"38",  x"a2",  x"06",  x"00", -- 3E50
         x"0d",  x"0c",  x"12",  x"23",  x"13",  x"18",  x"c7",  x"e1", -- 3E58
         x"04",  x"7e",  x"fe",  x"41",  x"38",  x"f4",  x"3e",  x"80", -- 3E60
         x"12",  x"c9",  x"04",  x"e1",  x"e5",  x"cd",  x"e3",  x"04", -- 3E68
         x"30",  x"fb",  x"28",  x"1b",  x"0f",  x"4f",  x"7e",  x"fe", -- 3E70
         x"61",  x"38",  x"06",  x"fe",  x"7b",  x"30",  x"02",  x"d6", -- 3E78
         x"20",  x"b9",  x"20",  x"e6",  x"23",  x"cd",  x"e3",  x"04", -- 3E80
         x"30",  x"ea",  x"2b",  x"f1",  x"78",  x"a7",  x"c9",  x"e1", -- 3E88
         x"7e",  x"c9",  x"1b",  x"13",  x"21",  x"00",  x"00",  x"1a", -- 3E90
         x"fe",  x"20",  x"28",  x"f7",  x"fe",  x"2d",  x"28",  x"13", -- 3E98
         x"d6",  x"30",  x"fe",  x"0a",  x"d0",  x"44",  x"4d",  x"29", -- 3EA0
         x"29",  x"09",  x"29",  x"06",  x"00",  x"4f",  x"09",  x"13", -- 3EA8
         x"1a",  x"18",  x"ed",  x"cd",  x"af",  x"de",  x"eb",  x"a7", -- 3EB0
         x"ed",  x"62",  x"ed",  x"52",  x"c9",  x"cd",  x"f5",  x"04", -- 3EB8
         x"fd",  x"e1",  x"cd",  x"41",  x"c6",  x"fd",  x"e5",  x"18", -- 3EC0
         x"35",  x"cd",  x"f5",  x"04",  x"ed",  x"b0",  x"18",  x"2e", -- 3EC8
         x"cd",  x"f5",  x"04",  x"cd",  x"3a",  x"cd",  x"18",  x"26", -- 3ED0
         x"cd",  x"f5",  x"04",  x"cd",  x"ae",  x"d6",  x"18",  x"03", -- 3ED8
         x"cd",  x"f5",  x"04",  x"cd",  x"34",  x"d8",  x"18",  x"16", -- 3EE0
         x"cd",  x"f5",  x"04",  x"cd",  x"8a",  x"d1",  x"18",  x"0e", -- 3EE8
         x"cd",  x"f5",  x"04",  x"cd",  x"cc",  x"d1",  x"18",  x"06", -- 3EF0
         x"cd",  x"f5",  x"04",  x"1a",  x"13",  x"87",  x"f5",  x"3a", -- 3EF8
         x"0e",  x"0a",  x"d3",  x"88",  x"dd",  x"cb",  x"04",  x"af", -- 3F00
         x"18",  x"05",  x"f5",  x"dd",  x"cb",  x"04",  x"ef",  x"d3", -- 3F08
         x"86",  x"f1",  x"c9",  x"02",  x"fe",  x"0d",  x"c4",  x"03", -- 3F10
         x"f0",  x"00",  x"fe",  x"20",  x"d0",  x"cd",  x"e9",  x"04", -- 3F18
         x"cd",  x"e9",  x"dd",  x"c3",  x"d7",  x"dd",  x"f5",  x"d5", -- 3F20
         x"db",  x"88",  x"5f",  x"f6",  x"85",  x"d3",  x"88",  x"dd", -- 3F28
         x"7e",  x"04",  x"57",  x"f6",  x"40",  x"e6",  x"5f",  x"dd", -- 3F30
         x"77",  x"04",  x"d3",  x"86",  x"cd",  x"fa",  x"db",  x"7a", -- 3F38
         x"dd",  x"77",  x"04",  x"d3",  x"86",  x"7b",  x"d3",  x"88", -- 3F40
         x"d1",  x"dc",  x"00",  x"00",  x"f1",  x"c9",  x"3a",  x"11", -- 3F48
         x"e0",  x"fe",  x"7f",  x"cc",  x"2f",  x"e0",  x"db",  x"88", -- 3F50
         x"e6",  x"fb",  x"0f",  x"17",  x"17",  x"0f",  x"d3",  x"88", -- 3F58
         x"cd",  x"4f",  x"c6",  x"c3",  x"54",  x"c8",  x"7f",  x"7f", -- 3F60
         x"42",  x"53",  x"41",  x"56",  x"45",  x"01",  x"3a",  x"80", -- 3F68
         x"b7",  x"32",  x"b1",  x"aa",  x"21",  x"a9",  x"d9",  x"e5", -- 3F70
         x"3a",  x"00",  x"03",  x"fe",  x"c3",  x"20",  x"14",  x"3a", -- 3F78
         x"03",  x"03",  x"fe",  x"c3",  x"20",  x"0d",  x"21",  x"5f", -- 3F80
         x"03",  x"5e",  x"23",  x"56",  x"21",  x"00",  x"04",  x"ed", -- 3F88
         x"52",  x"38",  x"18",  x"cd",  x"03",  x"f0",  x"23",  x"42", -- 3F90
         x"41",  x"53",  x"49",  x"43",  x"2d",  x"50",  x"72",  x"6f", -- 3F98
         x"67",  x"72",  x"61",  x"6d",  x"6d",  x"3f",  x"07",  x"0d", -- 3FA0
         x"0a",  x"00",  x"c9",  x"2a",  x"d7",  x"03",  x"7c",  x"e6", -- 3FA8
         x"80",  x"20",  x"e0",  x"22",  x"84",  x"b7",  x"cd",  x"03", -- 3FB0
         x"f0",  x"23",  x"0b",  x"25",  x"42",  x"53",  x"41",  x"56", -- 3FB8
         x"45",  x"20",  x"30",  x"33",  x"30",  x"30",  x"20",  x"00", -- 3FC0
         x"11",  x"70",  x"03",  x"ed",  x"53",  x"86",  x"b7",  x"cd", -- 3FC8
         x"03",  x"f0",  x"1b",  x"cd",  x"57",  x"d2",  x"21",  x"4e", -- 3FD0
         x"df",  x"01",  x"18",  x"00",  x"ed",  x"b0",  x"21",  x"f8", -- 3FD8
         x"df",  x"cd",  x"23",  x"cf",  x"d8",  x"cd",  x"57",  x"d2", -- 3FE0
         x"21",  x"00",  x"03",  x"22",  x"82",  x"b7",  x"7c",  x"32", -- 3FE8
         x"81",  x"b7",  x"eb",  x"cd",  x"03",  x"f0",  x"36",  x"c9", -- 3FF0
         x"4b",  x"43",  x"42",  x"00",  x"ff",  x"ff",  x"ff",  x"ff", -- 3FF8
         x"0c",  x"c0",  x"18",  x"1a",  x"c0",  x"46",  x"28",  x"c0", -- 4000
         x"42",  x"36",  x"c0",  x"40",  x"54",  x"6f",  x"70",  x"20", -- 4008
         x"6f",  x"66",  x"20",  x"54",  x"65",  x"78",  x"74",  x"3a", -- 4010
         x"20",  x"00",  x"45",  x"6e",  x"64",  x"20",  x"6f",  x"66", -- 4018
         x"20",  x"54",  x"65",  x"78",  x"74",  x"3a",  x"20",  x"00", -- 4020
         x"53",  x"74",  x"61",  x"72",  x"74",  x"20",  x"6f",  x"66", -- 4028
         x"20",  x"4d",  x"43",  x"3a",  x"20",  x"00",  x"41",  x"53", -- 4030
         x"4d",  x"2d",  x"4f",  x"66",  x"66",  x"73",  x"65",  x"74", -- 4038
         x"20",  x"3a",  x"20",  x"00",  x"f5",  x"db",  x"88",  x"e6", -- 4040
         x"5b",  x"d3",  x"88",  x"f1",  x"c9",  x"cd",  x"5a",  x"00", -- 4048
         x"ed",  x"b0",  x"18",  x"2c",  x"cd",  x"5a",  x"00",  x"ed", -- 4050
         x"b8",  x"18",  x"25",  x"cd",  x"5a",  x"00",  x"ed",  x"b1", -- 4058
         x"18",  x"1e",  x"cd",  x"5a",  x"00",  x"ed",  x"b9",  x"18", -- 4060
         x"17",  x"cd",  x"5a",  x"00",  x"be",  x"18",  x"11",  x"00", -- 4068
         x"cd",  x"5a",  x"00",  x"7e",  x"18",  x"0a",  x"cd",  x"5a", -- 4070
         x"00",  x"1a",  x"18",  x"04",  x"cd",  x"5a",  x"00",  x"77", -- 4078
         x"f5",  x"db",  x"88",  x"f6",  x"a4",  x"d3",  x"88",  x"f1", -- 4080
         x"c9",  x"06",  x"08",  x"0e",  x"80",  x"ed",  x"78",  x"fe", -- 4088
         x"f6",  x"28",  x"09",  x"fe",  x"f4",  x"28",  x"05",  x"04", -- 4090
         x"20",  x"f1",  x"18",  x"09",  x"16",  x"c3",  x"68",  x"3e", -- 4098
         x"02",  x"cd",  x"03",  x"f0",  x"26",  x"21",  x"44",  x"c0", -- 40A0
         x"11",  x"5a",  x"00",  x"01",  x"45",  x"00",  x"ed",  x"b0", -- 40A8
         x"c9",  x"7f",  x"7f",  x"41",  x"53",  x"4d",  x"1f",  x"cd", -- 40B0
         x"03",  x"f0",  x"23",  x"0c",  x"0a",  x"0a",  x"3e",  x"3e", -- 40B8
         x"20",  x"43",  x"41",  x"4f",  x"53",  x"2d",  x"41",  x"73", -- 40C0
         x"73",  x"65",  x"6d",  x"62",  x"6c",  x"65",  x"72",  x"20", -- 40C8
         x"32",  x"2e",  x"30",  x"20",  x"20",  x"60",  x"20",  x"4d", -- 40D0
         x"4c",  x"20",  x"31",  x"39",  x"39",  x"37",  x"2d",  x"32", -- 40D8
         x"30",  x"31",  x"38",  x"20",  x"3c",  x"3c",  x"00",  x"cd", -- 40E0
         x"89",  x"c0",  x"21",  x"08",  x"28",  x"22",  x"10",  x"00", -- 40E8
         x"21",  x"00",  x"02",  x"22",  x"18",  x"00",  x"22",  x"42", -- 40F0
         x"00",  x"24",  x"7c",  x"fe",  x"e0",  x"28",  x"13",  x"cd", -- 40F8
         x"86",  x"00",  x"4f",  x"2f",  x"cd",  x"92",  x"00",  x"cd", -- 4100
         x"86",  x"00",  x"2f",  x"b9",  x"79",  x"cd",  x"92",  x"00", -- 4108
         x"28",  x"e7",  x"22",  x"44",  x"00",  x"22",  x"46",  x"00", -- 4110
         x"26",  x"00",  x"22",  x"40",  x"00",  x"cd",  x"80",  x"c0", -- 4118
         x"cd",  x"fb",  x"c2",  x"3e",  x"06",  x"32",  x"a1",  x"b7", -- 4120
         x"11",  x"00",  x"c0",  x"06",  x"04",  x"1a",  x"13",  x"6f", -- 4128
         x"1a",  x"13",  x"67",  x"cd",  x"03",  x"f0",  x"45",  x"1a", -- 4130
         x"13",  x"6f",  x"26",  x"00",  x"7e",  x"23",  x"66",  x"6f", -- 4138
         x"cd",  x"03",  x"f0",  x"1a",  x"cd",  x"03",  x"f0",  x"2c", -- 4140
         x"10",  x"e3",  x"21",  x"0d",  x"06",  x"22",  x"9c",  x"b7", -- 4148
         x"21",  x"04",  x"04",  x"22",  x"9e",  x"b7",  x"3e",  x"11", -- 4150
         x"cd",  x"03",  x"f0",  x"00",  x"21",  x"00",  x"00",  x"22", -- 4158
         x"a0",  x"b7",  x"cd",  x"03",  x"f0",  x"17",  x"11",  x"00", -- 4160
         x"00",  x"d5",  x"cd",  x"03",  x"f0",  x"32",  x"eb",  x"cd", -- 4168
         x"03",  x"f0",  x"18",  x"d1",  x"38",  x"aa",  x"21",  x"82", -- 4170
         x"b7",  x"7a",  x"87",  x"85",  x"6f",  x"ed",  x"4b",  x"97", -- 4178
         x"b7",  x"71",  x"2c",  x"70",  x"14",  x"7a",  x"fe",  x"04", -- 4180
         x"20",  x"df",  x"2a",  x"86",  x"b7",  x"22",  x"42",  x"00", -- 4188
         x"2a",  x"88",  x"b7",  x"22",  x"40",  x"00",  x"2a",  x"82", -- 4190
         x"b7",  x"01",  x"00",  x"02",  x"a7",  x"ed",  x"42",  x"da", -- 4198
         x"20",  x"c1",  x"2a",  x"44",  x"00",  x"ed",  x"5b",  x"84", -- 41A0
         x"b7",  x"ed",  x"52",  x"38",  x"f2",  x"2a",  x"82",  x"b7", -- 41A8
         x"eb",  x"ed",  x"52",  x"38",  x"ea",  x"ed",  x"42",  x"38", -- 41B0
         x"e6",  x"eb",  x"3e",  x"0d",  x"cd",  x"92",  x"00",  x"23", -- 41B8
         x"22",  x"18",  x"00",  x"22",  x"1c",  x"00",  x"2a",  x"84", -- 41C0
         x"b7",  x"22",  x"44",  x"00",  x"cd",  x"23",  x"c4",  x"ed", -- 41C8
         x"62",  x"22",  x"20",  x"00",  x"cd",  x"dd",  x"c6",  x"cd", -- 41D0
         x"ce",  x"c4",  x"18",  x"0b",  x"7f",  x"7f",  x"52",  x"45", -- 41D8
         x"41",  x"53",  x"4d",  x"1f",  x"cd",  x"89",  x"c0",  x"af", -- 41E0
         x"32",  x"22",  x"00",  x"01",  x"f1",  x"83",  x"ed",  x"79", -- 41E8
         x"67",  x"6f",  x"06",  x"ff",  x"7e",  x"23",  x"fe",  x"7f", -- 41F0
         x"28",  x"04",  x"fe",  x"dd",  x"20",  x"05",  x"be",  x"20", -- 41F8
         x"02",  x"36",  x"00",  x"10",  x"ef",  x"cd",  x"fb",  x"c2", -- 4200
         x"3e",  x"0c",  x"cd",  x"03",  x"f0",  x"00",  x"21",  x"a2", -- 4208
         x"b7",  x"cb",  x"ce",  x"21",  x"3e",  x"00",  x"36",  x"40", -- 4210
         x"01",  x"80",  x"fc",  x"ed",  x"78",  x"fe",  x"a7",  x"20", -- 4218
         x"0d",  x"34",  x"01",  x"f1",  x"83",  x"ed",  x"78",  x"3c", -- 4220
         x"fe",  x"21",  x"38",  x"02",  x"cb",  x"ce",  x"01",  x"9e", -- 4228
         x"0d",  x"18",  x"0b",  x"dd",  x"dd",  x"4d",  x"45",  x"4e", -- 4230
         x"55",  x"1f",  x"e1",  x"01",  x"00",  x"26",  x"c5",  x"cd", -- 4238
         x"fb",  x"c2",  x"cd",  x"03",  x"f0",  x"23",  x"0c",  x"0a", -- 4240
         x"0a",  x"00",  x"06",  x"28",  x"cd",  x"03",  x"f0",  x"23", -- 4248
         x"5f",  x"00",  x"10",  x"f8",  x"cd",  x"28",  x"c3",  x"cd", -- 4250
         x"ad",  x"c3",  x"cd",  x"75",  x"c3",  x"3e",  x"1c",  x"32", -- 4258
         x"9f",  x"b7",  x"cd",  x"03",  x"f0",  x"2d",  x"21",  x"00", -- 4260
         x"ba",  x"c1",  x"cd",  x"03",  x"f0",  x"23",  x"02",  x"2a", -- 4268
         x"00",  x"cd",  x"03",  x"f0",  x"2a",  x"38",  x"4b",  x"3e", -- 4270
         x"dd",  x"ed",  x"b1",  x"e2",  x"c2",  x"c2",  x"ed",  x"a1", -- 4278
         x"20",  x"f7",  x"7e",  x"fe",  x"20",  x"38",  x"0f",  x"fe", -- 4280
         x"30",  x"38",  x"df",  x"fe",  x"5f",  x"30",  x"db",  x"cd", -- 4288
         x"55",  x"c5",  x"23",  x"0b",  x"18",  x"ec",  x"cd",  x"50", -- 4290
         x"c5",  x"18",  x"cf",  x"e1",  x"cd",  x"03",  x"f0",  x"19", -- 4298
         x"18",  x"06",  x"3e",  x"0b",  x"cd",  x"03",  x"f0",  x"00", -- 42A0
         x"3e",  x"02",  x"cd",  x"03",  x"f0",  x"00",  x"cd",  x"03", -- 42A8
         x"f0",  x"20",  x"cd",  x"28",  x"c3",  x"cd",  x"75",  x"c3", -- 42B0
         x"cd",  x"ad",  x"c3",  x"cd",  x"03",  x"f0",  x"23",  x"0d", -- 42B8
         x"2a",  x"00",  x"cd",  x"03",  x"f0",  x"17",  x"38",  x"da", -- 42C0
         x"13",  x"1a",  x"fe",  x"20",  x"28",  x"ed",  x"a7",  x"28", -- 42C8
         x"ea",  x"3e",  x"dd",  x"21",  x"00",  x"ba",  x"01",  x"00", -- 42D0
         x"26",  x"cd",  x"03",  x"f0",  x"1d",  x"30",  x"bd",  x"7e", -- 42D8
         x"23",  x"e5",  x"fe",  x"1f",  x"28",  x"10",  x"cd",  x"03", -- 42E0
         x"f0",  x"22",  x"38",  x"af",  x"21",  x"ae",  x"c2",  x"e3", -- 42E8
         x"e5",  x"cd",  x"03",  x"f0",  x"15",  x"c9",  x"21",  x"ae", -- 42F0
         x"c2",  x"e3",  x"e9",  x"21",  x"00",  x"00",  x"22",  x"9c", -- 42F8
         x"b7",  x"21",  x"28",  x"20",  x"18",  x"09",  x"21",  x"00", -- 4300
         x"01",  x"22",  x"9c",  x"b7",  x"21",  x"28",  x"1f",  x"22", -- 4308
         x"9e",  x"b7",  x"cd",  x"03",  x"f0",  x"20",  x"cd",  x"03", -- 4310
         x"f0",  x"23",  x"12",  x"00",  x"c9",  x"7e",  x"e6",  x"7f", -- 4318
         x"23",  x"cd",  x"03",  x"f0",  x"42",  x"10",  x"f6",  x"c9", -- 4320
         x"2a",  x"a0",  x"b7",  x"e5",  x"3e",  x"01",  x"32",  x"9d", -- 4328
         x"b7",  x"21",  x"01",  x"00",  x"22",  x"a0",  x"b7",  x"21", -- 4330
         x"f5",  x"b7",  x"7e",  x"fe",  x"21",  x"38",  x"1c",  x"cd", -- 4338
         x"03",  x"f0",  x"23",  x"41",  x"53",  x"4d",  x"3a",  x"20", -- 4340
         x"00",  x"06",  x"08",  x"cd",  x"1d",  x"c3",  x"3e",  x"2e", -- 4348
         x"cd",  x"03",  x"f0",  x"00",  x"06",  x"03",  x"cd",  x"1d", -- 4350
         x"c3",  x"18",  x"48",  x"cd",  x"03",  x"f0",  x"23",  x"3e", -- 4358
         x"3e",  x"20",  x"4b",  x"43",  x"2d",  x"41",  x"53",  x"4d", -- 4360
         x"20",  x"32",  x"2e",  x"30",  x"20",  x"3c",  x"3c",  x"20", -- 4368
         x"0d",  x"0a",  x"00",  x"18",  x"2e",  x"2a",  x"a0",  x"b7", -- 4370
         x"e5",  x"3e",  x"01",  x"32",  x"9d",  x"b7",  x"21",  x"1d", -- 4378
         x"00",  x"22",  x"a0",  x"b7",  x"cd",  x"03",  x"f0",  x"23", -- 4380
         x"46",  x"72",  x"65",  x"69",  x"3a",  x"00",  x"2a",  x"1e", -- 4388
         x"00",  x"ed",  x"5b",  x"1c",  x"00",  x"af",  x"ed",  x"52", -- 4390
         x"cd",  x"03",  x"f0",  x"1a",  x"cd",  x"03",  x"f0",  x"23", -- 4398
         x"08",  x"48",  x"00",  x"3e",  x"04",  x"32",  x"9d",  x"b7", -- 43A0
         x"e1",  x"22",  x"a0",  x"b7",  x"c9",  x"2a",  x"a0",  x"b7", -- 43A8
         x"e5",  x"3e",  x"01",  x"32",  x"9d",  x"b7",  x"21",  x"13", -- 43B0
         x"00",  x"22",  x"a0",  x"b7",  x"3e",  x"28",  x"cd",  x"03", -- 43B8
         x"f0",  x"00",  x"06",  x"09",  x"cd",  x"03",  x"f0",  x"2b", -- 43C0
         x"10",  x"fa",  x"3e",  x"14",  x"32",  x"a0",  x"b7",  x"3e", -- 43C8
         x"fe",  x"cd",  x"03",  x"f0",  x"49",  x"11",  x"14",  x"00", -- 43D0
         x"cd",  x"03",  x"f0",  x"32",  x"11",  x"1f",  x"c4",  x"01", -- 43D8
         x"04",  x"00",  x"1a",  x"13",  x"ed",  x"a1",  x"20",  x"2f", -- 43E0
         x"ea",  x"e2",  x"c3",  x"21",  x"3e",  x"00",  x"cb",  x"4e", -- 43E8
         x"28",  x"25",  x"cd",  x"03",  x"f0",  x"23",  x"3a",  x"00", -- 43F0
         x"3e",  x"01",  x"01",  x"f1",  x"80",  x"ed",  x"79",  x"ed", -- 43F8
         x"78",  x"cb",  x"47",  x"20",  x"fa",  x"04",  x"ed",  x"78", -- 4400
         x"cd",  x"55",  x"c5",  x"04",  x"ed",  x"78",  x"c6",  x"90", -- 4408
         x"27",  x"ce",  x"40",  x"27",  x"cd",  x"55",  x"c5",  x"3e", -- 4410
         x"29",  x"cd",  x"03",  x"f0",  x"00",  x"18",  x"84",  x"44", -- 4418
         x"49",  x"53",  x"4b",  x"22",  x"46",  x"00",  x"2b",  x"22", -- 4420
         x"1a",  x"00",  x"22",  x"1e",  x"00",  x"3e",  x"03",  x"c3", -- 4428
         x"92",  x"00",  x"dd",  x"dd",  x"51",  x"55",  x"49",  x"54", -- 4430
         x"1f",  x"cd",  x"fb",  x"c2",  x"21",  x"a1",  x"b7",  x"7e", -- 4438
         x"c6",  x"04",  x"77",  x"23",  x"cb",  x"8e",  x"e1",  x"ed", -- 4440
         x"5b",  x"7f",  x"b7",  x"3e",  x"02",  x"6f",  x"1e",  x"26", -- 4448
         x"c3",  x"09",  x"f0",  x"dd",  x"dd",  x"43",  x"4c",  x"45", -- 4450
         x"41",  x"52",  x"1f",  x"2a",  x"1c",  x"00",  x"ed",  x"5b", -- 4458
         x"18",  x"00",  x"a7",  x"ed",  x"52",  x"44",  x"4d",  x"2a", -- 4460
         x"1a",  x"00",  x"ed",  x"5b",  x"1e",  x"00",  x"ed",  x"52", -- 4468
         x"09",  x"7c",  x"b5",  x"28",  x"2b",  x"cd",  x"03",  x"f0", -- 4470
         x"23",  x"0d",  x"44",  x"65",  x"6c",  x"65",  x"74",  x"65", -- 4478
         x"20",  x"54",  x"65",  x"78",  x"74",  x"00",  x"cd",  x"0d", -- 4480
         x"c8",  x"38",  x"15",  x"cd",  x"ce",  x"c4",  x"2a",  x"18", -- 4488
         x"00",  x"22",  x"1c",  x"00",  x"2a",  x"1a",  x"00",  x"22", -- 4490
         x"1e",  x"00",  x"cd",  x"75",  x"c3",  x"cd",  x"d9",  x"c4", -- 4498
         x"2a",  x"44",  x"00",  x"ed",  x"5b",  x"46",  x"00",  x"a7", -- 44A0
         x"ed",  x"52",  x"c8",  x"cd",  x"03",  x"f0",  x"23",  x"0d", -- 44A8
         x"44",  x"65",  x"6c",  x"65",  x"74",  x"65",  x"20",  x"4c", -- 44B0
         x"61",  x"62",  x"65",  x"6c",  x"73",  x"00",  x"cd",  x"0d", -- 44B8
         x"c8",  x"d8",  x"cd",  x"e9",  x"c8",  x"2a",  x"44",  x"00", -- 44C0
         x"cd",  x"23",  x"c4",  x"c3",  x"30",  x"c9",  x"21",  x"f5", -- 44C8
         x"b7",  x"06",  x"0b",  x"36",  x"20",  x"23",  x"10",  x"fb", -- 44D0
         x"c9",  x"11",  x"00",  x"00",  x"ed",  x"53",  x"20",  x"00", -- 44D8
         x"c9",  x"dd",  x"dd",  x"53",  x"41",  x"56",  x"45",  x"1f", -- 44E0
         x"cd",  x"30",  x"c9",  x"ed",  x"5b",  x"1e",  x"00",  x"2a", -- 44E8
         x"1a",  x"00",  x"af",  x"ed",  x"52",  x"c8",  x"cd",  x"88", -- 44F0
         x"c8",  x"d8",  x"cd",  x"50",  x"c5",  x"cd",  x"d5",  x"c8", -- 44F8
         x"21",  x"00",  x"00",  x"cd",  x"03",  x"f0",  x"08",  x"d8", -- 4500
         x"ed",  x"5b",  x"1e",  x"00",  x"21",  x"80",  x"b7",  x"45", -- 4508
         x"3e",  x"1a",  x"2d",  x"77",  x"20",  x"fc",  x"cd",  x"8c", -- 4510
         x"00",  x"13",  x"77",  x"fe",  x"03",  x"28",  x"03",  x"23", -- 4518
         x"10",  x"f4",  x"dd",  x"7e",  x"02",  x"cd",  x"03",  x"f0", -- 4520
         x"1c",  x"cd",  x"03",  x"f0",  x"23",  x"08",  x"08",  x"00", -- 4528
         x"cd",  x"03",  x"f0",  x"2a",  x"01",  x"a0",  x"00",  x"38", -- 4530
         x"10",  x"2a",  x"1a",  x"00",  x"ed",  x"52",  x"38",  x"09", -- 4538
         x"d5",  x"cd",  x"03",  x"f0",  x"01",  x"d1",  x"d8",  x"18", -- 4540
         x"c3",  x"cd",  x"03",  x"f0",  x"09",  x"d4",  x"1d",  x"c6", -- 4548
         x"cd",  x"03",  x"f0",  x"2c",  x"c9",  x"cd",  x"03",  x"f0", -- 4550
         x"24",  x"c9",  x"dd",  x"dd",  x"4c",  x"4f",  x"41",  x"44", -- 4558
         x"1f",  x"3e",  x"08",  x"cd",  x"03",  x"f0",  x"49",  x"28", -- 4560
         x"07",  x"cd",  x"88",  x"c8",  x"d8",  x"cd",  x"50",  x"c5", -- 4568
         x"cd",  x"d9",  x"c4",  x"21",  x"00",  x"b7",  x"dd",  x"75", -- 4570
         x"05",  x"dd",  x"74",  x"06",  x"dd",  x"cb",  x"07",  x"c6", -- 4578
         x"21",  x"00",  x"00",  x"cd",  x"03",  x"f0",  x"0a",  x"30", -- 4580
         x"01",  x"c9",  x"af",  x"cd",  x"29",  x"c6",  x"38",  x"76", -- 4588
         x"3e",  x"08",  x"cd",  x"03",  x"f0",  x"49",  x"20",  x"1c", -- 4590
         x"3e",  x"02",  x"cd",  x"55",  x"c5",  x"11",  x"00",  x"00", -- 4598
         x"21",  x"00",  x"b7",  x"01",  x"0b",  x"00",  x"7e",  x"fe", -- 45A0
         x"20",  x"d4",  x"55",  x"c5",  x"ed",  x"a0",  x"ea",  x"a6", -- 45A8
         x"c5",  x"cd",  x"50",  x"c5",  x"dd",  x"36",  x"03",  x"02", -- 45B0
         x"ed",  x"5b",  x"1c",  x"00",  x"2a",  x"1e",  x"00",  x"a7", -- 45B8
         x"ed",  x"52",  x"28",  x"53",  x"e5",  x"cd",  x"29",  x"c6", -- 45C0
         x"e1",  x"38",  x"25",  x"01",  x"80",  x"00",  x"ed",  x"42", -- 45C8
         x"30",  x"02",  x"09",  x"4d",  x"21",  x"00",  x"b7",  x"7e", -- 45D0
         x"fe",  x"03",  x"28",  x"14",  x"fe",  x"1a",  x"28",  x"10", -- 45D8
         x"7e",  x"23",  x"eb",  x"cd",  x"92",  x"00",  x"eb",  x"13", -- 45E0
         x"0d",  x"20",  x"ec",  x"dd",  x"34",  x"03",  x"18",  x"cc", -- 45E8
         x"2a",  x"1c",  x"00",  x"eb",  x"cd",  x"74",  x"c9",  x"2a", -- 45F0
         x"1a",  x"00",  x"2b",  x"3e",  x"0a",  x"cd",  x"92",  x"00", -- 45F8
         x"2b",  x"3e",  x"0d",  x"cd",  x"92",  x"00",  x"cd",  x"03", -- 4600
         x"f0",  x"0b",  x"cd",  x"50",  x"c5",  x"3a",  x"22",  x"00", -- 4608
         x"b7",  x"28",  x"0a",  x"cd",  x"ef",  x"c7",  x"c9",  x"3c", -- 4610
         x"32",  x"22",  x"00",  x"18",  x"d3",  x"21",  x"00",  x"00", -- 4618
         x"11",  x"f5",  x"b7",  x"01",  x"0b",  x"00",  x"ed",  x"b0", -- 4620
         x"c9",  x"2e",  x"04",  x"20",  x"06",  x"dd",  x"cb",  x"07", -- 4628
         x"fe",  x"18",  x"26",  x"cd",  x"03",  x"f0",  x"2a",  x"d8", -- 4630
         x"dd",  x"7e",  x"03",  x"fe",  x"02",  x"20",  x"15",  x"dd", -- 4638
         x"cb",  x"07",  x"7e",  x"28",  x"0f",  x"dd",  x"cb",  x"07", -- 4640
         x"be",  x"3a",  x"10",  x"b7",  x"a7",  x"28",  x"05",  x"dd", -- 4648
         x"35",  x"03",  x"18",  x"05",  x"cd",  x"03",  x"f0",  x"05", -- 4650
         x"d8",  x"3e",  x"01",  x"3d",  x"dd",  x"7e",  x"02",  x"f5", -- 4658
         x"dd",  x"be",  x"03",  x"28",  x"08",  x"3c",  x"20",  x"21", -- 4660
         x"7d",  x"fe",  x"04",  x"20",  x"1c",  x"f1",  x"38",  x"08", -- 4668
         x"f5",  x"3e",  x"02",  x"cd",  x"03",  x"f0",  x"00",  x"f1", -- 4670
         x"f5",  x"cd",  x"03",  x"f0",  x"1c",  x"f1",  x"38",  x"0f", -- 4678
         x"cd",  x"03",  x"f0",  x"23",  x"3e",  x"20",  x"00",  x"a7", -- 4680
         x"c9",  x"f1",  x"37",  x"2c",  x"2d",  x"18",  x"e9",  x"28", -- 4688
         x"0b",  x"cd",  x"03",  x"f0",  x"23",  x"2a",  x"08",  x"08", -- 4690
         x"08",  x"00",  x"18",  x"97",  x"67",  x"2d",  x"28",  x"0a", -- 4698
         x"cd",  x"03",  x"f0",  x"23",  x"3f",  x"20",  x"07",  x"00", -- 46A0
         x"18",  x"89",  x"cd",  x"03",  x"f0",  x"23",  x"21",  x"0a", -- 46A8
         x"0d",  x"00",  x"a7",  x"c9",  x"dd",  x"dd",  x"56",  x"45", -- 46B0
         x"52",  x"49",  x"46",  x"59",  x"1f",  x"cd",  x"03",  x"f0", -- 46B8
         x"11",  x"c9",  x"dd",  x"dd",  x"4b",  x"45",  x"59",  x"01", -- 46C0
         x"b7",  x"20",  x"05",  x"cd",  x"03",  x"f0",  x"3a",  x"c9", -- 46C8
         x"7d",  x"b7",  x"28",  x"09",  x"fe",  x"d5",  x"28",  x"0c", -- 46D0
         x"cd",  x"03",  x"f0",  x"39",  x"c9",  x"21",  x"02",  x"c7", -- 46D8
         x"06",  x"02",  x"18",  x"05",  x"21",  x"fe",  x"c6",  x"06", -- 46E0
         x"0b",  x"11",  x"00",  x"b9",  x"af",  x"12",  x"13",  x"ed", -- 46E8
         x"a0",  x"03",  x"10",  x"f9",  x"eb",  x"36",  x"00",  x"23", -- 46F0
         x"7d",  x"fe",  x"9c",  x"20",  x"f8",  x"c9",  x"5b",  x"5c", -- 46F8
         x"5d",  x"7e",  x"05",  x"06",  x"7b",  x"7c",  x"7d",  x"60", -- 4700
         x"7f",  x"dd",  x"dd",  x"41",  x"53",  x"4d",  x"1f",  x"cd", -- 4708
         x"03",  x"f0",  x"23",  x"4f",  x"70",  x"74",  x"69",  x"6f", -- 4710
         x"6e",  x"73",  x"28",  x"2b",  x"2c",  x"31",  x"2c",  x"32", -- 4718
         x"2c",  x"42",  x"2c",  x"4c",  x"2c",  x"4f",  x"2c",  x"50", -- 4720
         x"2c",  x"53",  x"29",  x"3f",  x"3a",  x"00",  x"01",  x"26", -- 4728
         x"1a",  x"cd",  x"35",  x"c8",  x"d8",  x"11",  x"8f",  x"c7", -- 4730
         x"06",  x"08",  x"e5",  x"c5",  x"1a",  x"13",  x"01",  x"0d", -- 4738
         x"00",  x"ed",  x"b1",  x"37",  x"28",  x"01",  x"3f",  x"21", -- 4740
         x"3f",  x"00",  x"cb",  x"16",  x"c1",  x"e1",  x"10",  x"ea", -- 4748
         x"cd",  x"50",  x"c5",  x"3a",  x"3f",  x"00",  x"e6",  x"88", -- 4750
         x"fe",  x"88",  x"c8",  x"cd",  x"d9",  x"c4",  x"cd",  x"e9", -- 4758
         x"c8",  x"21",  x"30",  x"c9",  x"e5",  x"cd",  x"50",  x"c5", -- 4760
         x"2a",  x"1c",  x"00",  x"3e",  x"03",  x"cd",  x"92",  x"00", -- 4768
         x"2a",  x"18",  x"00",  x"e5",  x"21",  x"3f",  x"00",  x"7e", -- 4770
         x"cb",  x"a6",  x"be",  x"2b",  x"cb",  x"9e",  x"28",  x"02", -- 4778
         x"cb",  x"de",  x"e6",  x"84",  x"20",  x"06",  x"2a",  x"44", -- 4780
         x"00",  x"cd",  x"23",  x"c4",  x"c3",  x"bb",  x"cc",  x"32", -- 4788
         x"4f",  x"42",  x"53",  x"31",  x"2b",  x"50",  x"4c",  x"dd", -- 4790
         x"dd",  x"45",  x"44",  x"49",  x"54",  x"1f",  x"21",  x"ab", -- 4798
         x"c7",  x"11",  x"e0",  x"bf",  x"d5",  x"01",  x"20",  x"00", -- 47A0
         x"ed",  x"b0",  x"c9",  x"21",  x"5a",  x"c5",  x"16",  x"f1", -- 47A8
         x"18",  x"10",  x"dd",  x"dd",  x"51",  x"55",  x"49",  x"54", -- 47B0
         x"20",  x"01",  x"21",  x"cb",  x"c7",  x"32",  x"e7",  x"bf", -- 47B8
         x"16",  x"e1",  x"e3",  x"3e",  x"02",  x"6f",  x"cd",  x"03", -- 47C0
         x"f0",  x"26",  x"c9",  x"cd",  x"a5",  x"c0",  x"c3",  x"2e", -- 47C8
         x"c2",  x"cd",  x"03",  x"f0",  x"0c",  x"d0",  x"fe",  x"03", -- 47D0
         x"37",  x"c8",  x"fe",  x"13",  x"37",  x"3f",  x"c0",  x"cd", -- 47D8
         x"e5",  x"c7",  x"d8",  x"18",  x"f5",  x"cd",  x"03",  x"f0", -- 47E0
         x"04",  x"fe",  x"03",  x"37",  x"c8",  x"3f",  x"c9",  x"cd", -- 47E8
         x"03",  x"f0",  x"23",  x"0d",  x"3e",  x"3e",  x"3e",  x"20", -- 47F0
         x"4e",  x"6f",  x"20",  x"4d",  x"65",  x"6d",  x"6f",  x"72", -- 47F8
         x"79",  x"20",  x"3c",  x"3c",  x"3c",  x"07",  x"0a",  x"00", -- 4800
         x"af",  x"32",  x"22",  x"00",  x"c9",  x"cd",  x"03",  x"f0", -- 4808
         x"23",  x"20",  x"28",  x"59",  x"2f",  x"4e",  x"29",  x"20", -- 4810
         x"3f",  x"20",  x"00",  x"cd",  x"e5",  x"c7",  x"38",  x"0c", -- 4818
         x"cd",  x"89",  x"d6",  x"fe",  x"59",  x"28",  x"05",  x"fe", -- 4820
         x"4e",  x"20",  x"f0",  x"37",  x"f5",  x"cd",  x"55",  x"c5", -- 4828
         x"cd",  x"50",  x"c5",  x"f1",  x"c9",  x"78",  x"32",  x"a0", -- 4830
         x"b7",  x"cd",  x"e5",  x"c7",  x"30",  x"05",  x"cd",  x"50", -- 4838
         x"c5",  x"37",  x"c9",  x"fe",  x"2e",  x"28",  x"1f",  x"fe", -- 4840
         x"05",  x"28",  x"20",  x"fe",  x"20",  x"30",  x"26",  x"fe", -- 4848
         x"08",  x"28",  x"22",  x"fe",  x"09",  x"28",  x"1e",  x"fe", -- 4850
         x"0d",  x"20",  x"de",  x"3a",  x"a1",  x"b7",  x"57",  x"58", -- 4858
         x"cd",  x"03",  x"f0",  x"32",  x"a7",  x"c9",  x"79",  x"fe", -- 4860
         x"10",  x"20",  x"08",  x"78",  x"c6",  x"08",  x"32",  x"a0", -- 4868
         x"b7",  x"18",  x"06",  x"3e",  x"2e",  x"cd",  x"03",  x"f0", -- 4870
         x"00",  x"21",  x"a0",  x"b7",  x"7e",  x"b8",  x"30",  x"01", -- 4878
         x"78",  x"b9",  x"38",  x"01",  x"79",  x"77",  x"18",  x"b1", -- 4880
         x"11",  x"cd",  x"c8",  x"cd",  x"03",  x"f0",  x"23",  x"0a", -- 4888
         x"0b",  x"4e",  x"61",  x"6d",  x"65",  x"20",  x"3a",  x"00", -- 4890
         x"7b",  x"a7",  x"0e",  x"11",  x"28",  x"13",  x"0d",  x"21", -- 4898
         x"f5",  x"b7",  x"06",  x"08",  x"7e",  x"23",  x"cd",  x"03", -- 48A0
         x"f0",  x"42",  x"10",  x"f8",  x"eb",  x"cd",  x"03",  x"f0", -- 48A8
         x"45",  x"06",  x"06",  x"d5",  x"cd",  x"35",  x"c8",  x"d1", -- 48B0
         x"d8",  x"7b",  x"a7",  x"28",  x"0a",  x"e5",  x"11",  x"00", -- 48B8
         x"00",  x"01",  x"0b",  x"00",  x"ed",  x"b0",  x"e1",  x"3e", -- 48C0
         x"13",  x"32",  x"a0",  x"b7",  x"c9",  x"41",  x"53",  x"4d", -- 48C8
         x"00",  x"4b",  x"43",  x"43",  x"00",  x"11",  x"80",  x"b7", -- 48D0
         x"af",  x"1d",  x"12",  x"20",  x"fc",  x"dd",  x"73",  x"05", -- 48D8
         x"dd",  x"72",  x"06",  x"01",  x"0b",  x"00",  x"ed",  x"b0", -- 48E0
         x"c9",  x"2a",  x"1a",  x"00",  x"ed",  x"4b",  x"1e",  x"00", -- 48E8
         x"af",  x"ed",  x"42",  x"44",  x"4d",  x"c8",  x"2a",  x"1e", -- 48F0
         x"00",  x"3e",  x"0d",  x"cd",  x"71",  x"00",  x"20",  x"10", -- 48F8
         x"1b",  x"e2",  x"10",  x"c9",  x"7a",  x"b3",  x"20",  x"f1", -- 4900
         x"cd",  x"86",  x"00",  x"fe",  x"0a",  x"20",  x"01",  x"23", -- 4908
         x"cd",  x"14",  x"c9",  x"c9",  x"ed",  x"5b",  x"1e",  x"00", -- 4910
         x"d5",  x"af",  x"ed",  x"52",  x"44",  x"4d",  x"e1",  x"ed", -- 4918
         x"5b",  x"1c",  x"00",  x"28",  x"03",  x"cd",  x"63",  x"00", -- 4920
         x"ed",  x"53",  x"1c",  x"00",  x"22",  x"1e",  x"00",  x"c9", -- 4928
         x"cd",  x"d9",  x"c4",  x"2a",  x"1c",  x"00",  x"ed",  x"4b", -- 4930
         x"18",  x"00",  x"af",  x"ed",  x"42",  x"44",  x"4d",  x"c8", -- 4938
         x"03",  x"2a",  x"1c",  x"00",  x"2b",  x"cd",  x"86",  x"00", -- 4940
         x"fe",  x"0a",  x"20",  x"02",  x"2b",  x"0b",  x"cd",  x"86", -- 4948
         x"00",  x"fe",  x"0d",  x"20",  x"02",  x"2b",  x"0b",  x"3e", -- 4950
         x"0d",  x"cd",  x"78",  x"00",  x"1b",  x"20",  x"08",  x"e2", -- 4958
         x"66",  x"c9",  x"7a",  x"b3",  x"20",  x"f1",  x"23",  x"23", -- 4960
         x"cd",  x"86",  x"00",  x"fe",  x"0a",  x"20",  x"01",  x"23", -- 4968
         x"eb",  x"2a",  x"1c",  x"00",  x"e5",  x"af",  x"ed",  x"52", -- 4970
         x"44",  x"4d",  x"e1",  x"ed",  x"5b",  x"1e",  x"00",  x"1b", -- 4978
         x"2b",  x"c4",  x"6a",  x"00",  x"13",  x"ed",  x"53",  x"1e", -- 4980
         x"00",  x"23",  x"22",  x"1c",  x"00",  x"c9",  x"dd",  x"dd", -- 4988
         x"48",  x"45",  x"4c",  x"50",  x"1f",  x"cd",  x"03",  x"f0", -- 4990
         x"23",  x"10",  x"02",  x"45",  x"72",  x"72",  x"6f",  x"72", -- 4998
         x"73",  x"3a",  x"0a",  x"02",  x"31",  x"2d",  x"53",  x"65", -- 49A0
         x"6d",  x"69",  x"6b",  x"6f",  x"6c",  x"6f",  x"6e",  x"3f", -- 49A8
         x"0a",  x"02",  x"32",  x"2d",  x"4d",  x"61",  x"72",  x"6b", -- 49B0
         x"65",  x"20",  x"32",  x"2a",  x"0a",  x"02",  x"33",  x"2d", -- 49B8
         x"4d",  x"61",  x"72",  x"6b",  x"65",  x"20",  x"66",  x"65", -- 49C0
         x"68",  x"6c",  x"74",  x"0a",  x"02",  x"34",  x"2d",  x"53", -- 49C8
         x"79",  x"6e",  x"74",  x"61",  x"78",  x"66",  x"65",  x"68", -- 49D0
         x"6c",  x"65",  x"72",  x"0a",  x"02",  x"35",  x"2d",  x"5a", -- 49D8
         x"61",  x"68",  x"6c",  x"65",  x"6e",  x"66",  x"6f",  x"72", -- 49E0
         x"6d",  x"61",  x"74",  x"3f",  x"0a",  x"02",  x"36",  x"2d", -- 49E8
         x"42",  x"65",  x"72",  x"65",  x"69",  x"63",  x"68",  x"20", -- 49F0
         x"76",  x"65",  x"72",  x"6c",  x"61",  x"73",  x"73",  x"65", -- 49F8
         x"6e",  x"0a",  x"02",  x"37",  x"2d",  x"45",  x"51",  x"55", -- 4A00
         x"20",  x"6f",  x"68",  x"6e",  x"65",  x"20",  x"4d",  x"61", -- 4A08
         x"72",  x"6b",  x"65",  x"0a",  x"02",  x"38",  x"2d",  x"5a", -- 4A10
         x"65",  x"69",  x"63",  x"68",  x"65",  x"6e",  x"6b",  x"65", -- 4A18
         x"74",  x"74",  x"65",  x"0a",  x"02",  x"39",  x"2d",  x"4f", -- 4A20
         x"70",  x"65",  x"72",  x"61",  x"6e",  x"64",  x"65",  x"6e", -- 4A28
         x"66",  x"65",  x"68",  x"6c",  x"65",  x"72",  x"0a",  x"02", -- 4A30
         x"41",  x"2d",  x"46",  x"6c",  x"61",  x"67",  x"73",  x"0a", -- 4A38
         x"02",  x"42",  x"2d",  x"52",  x"65",  x"63",  x"68",  x"65", -- 4A40
         x"6e",  x"7a",  x"65",  x"69",  x"63",  x"68",  x"65",  x"6e", -- 4A48
         x"0a",  x"02",  x"43",  x"2d",  x"44",  x"69",  x"76",  x"69", -- 4A50
         x"73",  x"69",  x"6f",  x"6e",  x"2f",  x"30",  x"0a",  x"02", -- 4A58
         x"44",  x"2d",  x"4d",  x"61",  x"72",  x"6b",  x"65",  x"20", -- 4A60
         x"64",  x"6f",  x"70",  x"70",  x"65",  x"6c",  x"74",  x"0a", -- 4A68
         x"02",  x"45",  x"2d",  x"49",  x"6e",  x"64",  x"65",  x"78", -- 4A70
         x"72",  x"65",  x"67",  x"69",  x"73",  x"74",  x"65",  x"72", -- 4A78
         x"0a",  x"02",  x"00",  x"c9",  x"dd",  x"dd",  x"4c",  x"41", -- 4A80
         x"42",  x"45",  x"4c",  x"1f",  x"1e",  x"00",  x"cd",  x"8b", -- 4A88
         x"c8",  x"d8",  x"11",  x"23",  x"00",  x"01",  x"08",  x"00", -- 4A90
         x"ed",  x"b0",  x"21",  x"23",  x"00",  x"cd",  x"5d",  x"d6", -- 4A98
         x"38",  x"06",  x"cd",  x"03",  x"f0",  x"1a",  x"18",  x"0e", -- 4AA0
         x"cd",  x"03",  x"f0",  x"23",  x"6e",  x"6f",  x"74",  x"20", -- 4AA8
         x"66",  x"6f",  x"75",  x"6e",  x"64",  x"00",  x"c3",  x"50", -- 4AB0
         x"c5",  x"dd",  x"dd",  x"4c",  x"42",  x"4c",  x"49",  x"53", -- 4AB8
         x"54",  x"01",  x"b7",  x"0e",  x"03",  x"28",  x"01",  x"4d", -- 4AC0
         x"2a",  x"46",  x"00",  x"c5",  x"eb",  x"2a",  x"44",  x"00", -- 4AC8
         x"37",  x"ed",  x"52",  x"38",  x"46",  x"eb",  x"cd",  x"86", -- 4AD0
         x"00",  x"5f",  x"23",  x"cd",  x"86",  x"00",  x"57",  x"23", -- 4AD8
         x"eb",  x"cd",  x"03",  x"f0",  x"1a",  x"cd",  x"8c",  x"00", -- 4AE0
         x"13",  x"3d",  x"20",  x"07",  x"cd",  x"03",  x"f0",  x"23", -- 4AE8
         x"08",  x"2a",  x"00",  x"eb",  x"06",  x"08",  x"cd",  x"86", -- 4AF0
         x"00",  x"23",  x"fe",  x"3a",  x"28",  x"0f",  x"cd",  x"55", -- 4AF8
         x"c5",  x"10",  x"f3",  x"cd",  x"86",  x"00",  x"23",  x"fe", -- 4B00
         x"3a",  x"20",  x"f8",  x"18",  x"06",  x"cd",  x"03",  x"f0", -- 4B08
         x"2b",  x"10",  x"fa",  x"cd",  x"d1",  x"c7",  x"38",  x"03", -- 4B10
         x"0d",  x"20",  x"b1",  x"c1",  x"f5",  x"cd",  x"50",  x"c5", -- 4B18
         x"f1",  x"30",  x"a8",  x"c9",  x"cd",  x"86",  x"00",  x"fe", -- 4B20
         x"20",  x"28",  x"03",  x"fe",  x"09",  x"c0",  x"23",  x"18", -- 4B28
         x"f3",  x"cd",  x"86",  x"00",  x"fe",  x"20",  x"30",  x"2b", -- 4B30
         x"23",  x"e5",  x"d5",  x"c5",  x"23",  x"13",  x"cd",  x"8c", -- 4B38
         x"00",  x"cd",  x"75",  x"d6",  x"38",  x"0c",  x"47",  x"cd", -- 4B40
         x"86",  x"00",  x"cd",  x"75",  x"d6",  x"b8",  x"20",  x"0f", -- 4B48
         x"18",  x"ea",  x"cd",  x"86",  x"00",  x"cd",  x"75",  x"d6", -- 4B50
         x"30",  x"05",  x"c1",  x"e1",  x"e1",  x"b7",  x"c9",  x"c1", -- 4B58
         x"d1",  x"e1",  x"2b",  x"37",  x"c9",  x"3a",  x"80",  x"a8", -- 4B60
         x"fe",  x"20",  x"28",  x"15",  x"3e",  x"2a",  x"32",  x"81", -- 4B68
         x"a8",  x"2a",  x"4e",  x"00",  x"7d",  x"c6",  x"01",  x"27", -- 4B70
         x"6f",  x"7c",  x"ce",  x"00",  x"27",  x"67",  x"22",  x"4e", -- 4B78
         x"00",  x"21",  x"80",  x"a8",  x"11",  x"00",  x"60",  x"3a", -- 4B80
         x"3f",  x"00",  x"e6",  x"20",  x"28",  x"02",  x"16",  x"27", -- 4B88
         x"7e",  x"23",  x"fe",  x"0d",  x"28",  x"07",  x"cd",  x"9a", -- 4B90
         x"d6",  x"7b",  x"ba",  x"38",  x"f3",  x"3e",  x"0d",  x"cd", -- 4B98
         x"9a",  x"d6",  x"21",  x"80",  x"a8",  x"06",  x"10",  x"36", -- 4BA0
         x"20",  x"23",  x"10",  x"fb",  x"36",  x"0d",  x"c9",  x"21", -- 4BA8
         x"82",  x"a8",  x"7a",  x"cd",  x"b7",  x"cb",  x"7b",  x"f5", -- 4BB0
         x"1f",  x"1f",  x"1f",  x"1f",  x"cd",  x"c0",  x"cb",  x"f1", -- 4BB8
         x"e6",  x"0f",  x"c6",  x"90",  x"27",  x"ce",  x"40",  x"27", -- 4BC0
         x"77",  x"23",  x"c9",  x"cd",  x"eb",  x"cc",  x"3a",  x"3e", -- 4BC8
         x"00",  x"cb",  x"57",  x"28",  x"04",  x"e1",  x"c3",  x"50", -- 4BD0
         x"c5",  x"3a",  x"3f",  x"00",  x"17",  x"30",  x"36",  x"e5", -- 4BD8
         x"f5",  x"1f",  x"1f",  x"dc",  x"65",  x"cb",  x"f1",  x"cb", -- 4BE0
         x"6f",  x"20",  x"08",  x"3a",  x"80",  x"a8",  x"fe",  x"20", -- 4BE8
         x"c4",  x"65",  x"cb",  x"cd",  x"a2",  x"cb",  x"ed",  x"5b", -- 4BF0
         x"4c",  x"00",  x"cd",  x"af",  x"cb",  x"23",  x"22",  x"48", -- 4BF8
         x"00",  x"e1",  x"e5",  x"11",  x"90",  x"a8",  x"06",  x"50", -- 4C00
         x"cd",  x"86",  x"00",  x"12",  x"fe",  x"0d",  x"28",  x"04", -- 4C08
         x"13",  x"23",  x"10",  x"f4",  x"e1",  x"cd",  x"03",  x"f0", -- 4C10
         x"2a",  x"30",  x"09",  x"3a",  x"3f",  x"00",  x"cb",  x"67", -- 4C18
         x"20",  x"75",  x"e1",  x"c9",  x"cd",  x"86",  x"00",  x"fe", -- 4C20
         x"03",  x"20",  x"a0",  x"cd",  x"a2",  x"cb",  x"21",  x"3f", -- 4C28
         x"00",  x"7e",  x"17",  x"30",  x"6e",  x"e6",  x"20",  x"20", -- 4C30
         x"5e",  x"cd",  x"03",  x"f0",  x"23",  x"0a",  x"45",  x"72", -- 4C38
         x"72",  x"6f",  x"72",  x"73",  x"3a",  x"20",  x"00",  x"2a", -- 4C40
         x"4e",  x"00",  x"cd",  x"03",  x"f0",  x"1a",  x"cd",  x"50", -- 4C48
         x"c5",  x"cd",  x"4f",  x"d6",  x"38",  x"14",  x"cd",  x"03", -- 4C50
         x"f0",  x"23",  x"53",  x"74",  x"61",  x"72",  x"74",  x"20", -- 4C58
         x"3a",  x"20",  x"00",  x"cd",  x"03",  x"f0",  x"1a",  x"cd", -- 4C60
         x"50",  x"c5",  x"cd",  x"03",  x"f0",  x"23",  x"45",  x"6e", -- 4C68
         x"64",  x"2b",  x"31",  x"20",  x"3a",  x"20",  x"00",  x"2a", -- 4C70
         x"4c",  x"00",  x"cd",  x"03",  x"f0",  x"1a",  x"cd",  x"50", -- 4C78
         x"c5",  x"2a",  x"4e",  x"00",  x"7c",  x"b5",  x"20",  x"19", -- 4C80
         x"21",  x"3e",  x"00",  x"cb",  x"5e",  x"28",  x"12",  x"23", -- 4C88
         x"36",  x"90",  x"cd",  x"d1",  x"d6",  x"18",  x"24",  x"01", -- 4C90
         x"a0",  x"00",  x"cd",  x"03",  x"f0",  x"09",  x"cd",  x"50", -- 4C98
         x"c5",  x"e1",  x"c9",  x"cb",  x"fe",  x"cd",  x"03",  x"f0", -- 4CA0
         x"23",  x"45",  x"6e",  x"64",  x"20",  x"50",  x"61",  x"73", -- 4CA8
         x"73",  x"20",  x"31",  x"0d",  x"0a",  x"0a",  x"00",  x"cb", -- 4CB0
         x"5e",  x"20",  x"af",  x"21",  x"3e",  x"00",  x"cb",  x"be", -- 4CB8
         x"cb",  x"96",  x"cd",  x"a2",  x"cb",  x"21",  x"00",  x"00", -- 4CC0
         x"22",  x"4e",  x"00",  x"22",  x"50",  x"00",  x"3a",  x"3f", -- 4CC8
         x"00",  x"e6",  x"82",  x"fe",  x"82",  x"20",  x"07",  x"21", -- 4CD0
         x"08",  x"f0",  x"cd",  x"03",  x"f0",  x"1e",  x"e1",  x"e5", -- 4CD8
         x"fd",  x"2a",  x"42",  x"00",  x"fd",  x"22",  x"4c",  x"00", -- 4CE0
         x"c3",  x"ce",  x"cb",  x"3a",  x"3e",  x"00",  x"a7",  x"fa", -- 4CE8
         x"68",  x"ce",  x"cd",  x"86",  x"00",  x"0e",  x"ff",  x"cd", -- 4CF0
         x"89",  x"d6",  x"30",  x"19",  x"cd",  x"24",  x"cb",  x"fe", -- 4CF8
         x"0d",  x"28",  x"0f",  x"fe",  x"3b",  x"28",  x"0b",  x"cd", -- 4D00
         x"89",  x"d6",  x"d2",  x"a6",  x"cd",  x"3e",  x"31",  x"32", -- 4D08
         x"80",  x"a8",  x"c3",  x"68",  x"ce",  x"0c",  x"54",  x"5d", -- 4D10
         x"cd",  x"39",  x"cb",  x"eb",  x"fe",  x"3a",  x"20",  x"06", -- 4D18
         x"23",  x"cd",  x"86",  x"00",  x"18",  x"f6",  x"e5",  x"d5", -- 4D20
         x"a7",  x"ed",  x"52",  x"23",  x"23",  x"23",  x"e5",  x"2a", -- 4D28
         x"1e",  x"00",  x"ed",  x"5b",  x"1c",  x"00",  x"ed",  x"52", -- 4D30
         x"d1",  x"37",  x"ed",  x"52",  x"e1",  x"30",  x"0c",  x"cd", -- 4D38
         x"ef",  x"c7",  x"21",  x"3e",  x"00",  x"cb",  x"d6",  x"e1", -- 4D40
         x"c3",  x"68",  x"ce",  x"c5",  x"cd",  x"2d",  x"d6",  x"c1", -- 4D48
         x"d1",  x"38",  x"1c",  x"2b",  x"3a",  x"3f",  x"00",  x"17", -- 4D50
         x"30",  x"0d",  x"cd",  x"86",  x"00",  x"3d",  x"20",  x"0c", -- 4D58
         x"3e",  x"44",  x"32",  x"80",  x"a8",  x"18",  x"05",  x"3e", -- 4D60
         x"01",  x"cd",  x"92",  x"00",  x"eb",  x"18",  x"8d",  x"3a", -- 4D68
         x"3f",  x"00",  x"17",  x"38",  x"f7",  x"d5",  x"3e",  x"3a", -- 4D70
         x"cd",  x"92",  x"00",  x"2b",  x"1b",  x"cd",  x"8c",  x"00", -- 4D78
         x"fe",  x"3a",  x"28",  x"f8",  x"cd",  x"89",  x"d6",  x"cd", -- 4D80
         x"92",  x"00",  x"2b",  x"fe",  x"20",  x"30",  x"ed",  x"ed", -- 4D88
         x"5b",  x"4c",  x"00",  x"7a",  x"cd",  x"92",  x"00",  x"2b", -- 4D90
         x"7b",  x"cd",  x"92",  x"00",  x"cd",  x"23",  x"c4",  x"cd", -- 4D98
         x"75",  x"c3",  x"e1",  x"c3",  x"fc",  x"cc",  x"11",  x"00", -- 4DA0
         x"00",  x"d6",  x"40",  x"47",  x"83",  x"5f",  x"7a",  x"82", -- 4DA8
         x"80",  x"57",  x"23",  x"cd",  x"86",  x"00",  x"cd",  x"89", -- 4DB0
         x"d6",  x"30",  x"ee",  x"e5",  x"fe",  x"20",  x"28",  x"0c", -- 4DB8
         x"fe",  x"09",  x"28",  x"08",  x"fe",  x"3b",  x"28",  x"04", -- 4DC0
         x"fe",  x"0d",  x"20",  x"60",  x"a7",  x"21",  x"2b",  x"4b", -- 4DC8
         x"ed",  x"52",  x"28",  x"18",  x"7a",  x"01",  x"28",  x"00", -- 4DD0
         x"21",  x"cf",  x"d5",  x"ed",  x"b1",  x"20",  x"33",  x"3e", -- 4DD8
         x"06",  x"b9",  x"38",  x"28",  x"7a",  x"83",  x"fe",  x"73", -- 4DE0
         x"38",  x"fb",  x"18",  x"e9",  x"79",  x"b7",  x"3e",  x"37", -- 4DE8
         x"20",  x"3c",  x"e1",  x"cd",  x"d2",  x"d2",  x"3a",  x"3f", -- 4DF0
         x"00",  x"17",  x"38",  x"6c",  x"e5",  x"2a",  x"46",  x"00", -- 4DF8
         x"7b",  x"cd",  x"92",  x"00",  x"23",  x"7a",  x"cd",  x"92", -- 4E00
         x"00",  x"e1",  x"18",  x"5c",  x"01",  x"27",  x"00",  x"09", -- 4E08
         x"53",  x"5e",  x"7a",  x"16",  x"00",  x"21",  x"31",  x"d5", -- 4E10
         x"19",  x"46",  x"21",  x"80",  x"d5",  x"19",  x"4e",  x"e6", -- 4E18
         x"07",  x"57",  x"79",  x"0f",  x"0f",  x"0f",  x"0f",  x"e6", -- 4E20
         x"07",  x"92",  x"28",  x"05",  x"3e",  x"34",  x"32",  x"80", -- 4E28
         x"a8",  x"e1",  x"20",  x"34",  x"c5",  x"af",  x"32",  x"4a", -- 4E30
         x"00",  x"79",  x"e6",  x"0f",  x"fe",  x"0d",  x"28",  x"1d", -- 4E38
         x"fe",  x"0e",  x"28",  x"19",  x"e5",  x"cd",  x"87",  x"d2", -- 4E40
         x"dc",  x"0f",  x"d2",  x"2b",  x"cd",  x"86",  x"00",  x"23", -- 4E48
         x"fe",  x"2c",  x"cc",  x"0f",  x"d2",  x"3a",  x"4a",  x"00", -- 4E50
         x"b7",  x"c4",  x"50",  x"d2",  x"e1",  x"f1",  x"f5",  x"3e", -- 4E58
         x"ed",  x"fc",  x"50",  x"d2",  x"c1",  x"cd",  x"7f",  x"ce", -- 4E60
         x"fd",  x"22",  x"4c",  x"00",  x"3e",  x"0d",  x"c5",  x"01", -- 4E68
         x"00",  x"01",  x"cd",  x"71",  x"00",  x"cd",  x"86",  x"00", -- 4E70
         x"fe",  x"0a",  x"20",  x"01",  x"23",  x"c1",  x"c9",  x"e5", -- 4E78
         x"c5",  x"3e",  x"0f",  x"a1",  x"21",  x"99",  x"ce",  x"11", -- 4E80
         x"f3",  x"d4",  x"3c",  x"06",  x"00",  x"f5",  x"1a",  x"13", -- 4E88
         x"4f",  x"09",  x"f1",  x"3d",  x"20",  x"f7",  x"c1",  x"e3", -- 4E90
         x"c9",  x"3a",  x"3e",  x"00",  x"cb",  x"ff",  x"32",  x"3e", -- 4E98
         x"00",  x"c9",  x"3e",  x"cb",  x"cd",  x"50",  x"d2",  x"cd", -- 4EA0
         x"0f",  x"d2",  x"7b",  x"fe",  x"08",  x"d2",  x"7a",  x"d0", -- 4EA8
         x"07",  x"07",  x"07",  x"80",  x"47",  x"cd",  x"0f",  x"d2", -- 4EB0
         x"28",  x"2b",  x"4f",  x"cd",  x"2d",  x"d2",  x"30",  x"2a", -- 4EB8
         x"3e",  x"06",  x"b9",  x"20",  x"20",  x"78",  x"e6",  x"c0", -- 4EC0
         x"fe",  x"40",  x"28",  x"1e",  x"2b",  x"cd",  x"86",  x"00", -- 4EC8
         x"23",  x"fe",  x"2c",  x"20",  x"15",  x"cd",  x"0f",  x"d2", -- 4ED0
         x"28",  x"0b",  x"fe",  x"06",  x"28",  x"07",  x"4f",  x"3a", -- 4ED8
         x"54",  x"00",  x"a7",  x"28",  x"05",  x"3e",  x"45",  x"32", -- 4EE0
         x"80",  x"a8",  x"79",  x"c3",  x"44",  x"d2",  x"3a",  x"54", -- 4EE8
         x"00",  x"90",  x"c8",  x"e6",  x"0f",  x"28",  x"0b",  x"79", -- 4EF0
         x"ab",  x"e6",  x"04",  x"c0",  x"3e",  x"07",  x"b9",  x"c8", -- 4EF8
         x"bb",  x"c8",  x"3e",  x"45",  x"c3",  x"e3",  x"d1",  x"3e", -- 4F00
         x"06",  x"b9",  x"c0",  x"bb",  x"c0",  x"3e",  x"39",  x"18", -- 4F08
         x"f3",  x"e5",  x"af",  x"32",  x"4a",  x"00",  x"cd",  x"0f", -- 4F10
         x"d2",  x"28",  x"31",  x"4f",  x"3a",  x"54",  x"00",  x"47", -- 4F18
         x"cd",  x"0f",  x"d2",  x"28",  x"5d",  x"5f",  x"81",  x"fe", -- 4F20
         x"0f",  x"d2",  x"f0",  x"cf",  x"e1",  x"7b",  x"c6",  x"40", -- 4F28
         x"c5",  x"47",  x"79",  x"cd",  x"41",  x"d2",  x"c1",  x"cd", -- 4F30
         x"07",  x"cf",  x"3a",  x"4a",  x"00",  x"b7",  x"c8",  x"3e", -- 4F38
         x"06",  x"bb",  x"28",  x"03",  x"b9",  x"20",  x"a7",  x"3a", -- 4F40
         x"4b",  x"00",  x"18",  x"47",  x"d1",  x"3a",  x"59",  x"00", -- 4F48
         x"3c",  x"28",  x"03",  x"3c",  x"18",  x"3d",  x"ed",  x"4b", -- 4F50
         x"52",  x"00",  x"cd",  x"0f",  x"d2",  x"ed",  x"43",  x"52", -- 4F58
         x"00",  x"fe",  x"07",  x"20",  x"07",  x"3e",  x"32",  x"cd", -- 4F60
         x"50",  x"d2",  x"18",  x"43",  x"fe",  x"20",  x"06",  x"22", -- 4F68
         x"28",  x"0a",  x"f5",  x"3e",  x"ed",  x"cd",  x"50",  x"d2", -- 4F70
         x"f1",  x"c6",  x"43",  x"47",  x"78",  x"cd",  x"50",  x"d2", -- 4F78
         x"18",  x"2d",  x"e1",  x"fe",  x"28",  x"20",  x"0f",  x"32", -- 4F80
         x"4a",  x"00",  x"3a",  x"59",  x"00",  x"fe",  x"ff",  x"28", -- 4F88
         x"05",  x"c6",  x"0a",  x"c3",  x"50",  x"d2",  x"cd",  x"d2", -- 4F90
         x"d2",  x"3a",  x"59",  x"00",  x"fe",  x"07",  x"20",  x"12", -- 4F98
         x"3a",  x"4a",  x"00",  x"fe",  x"28",  x"20",  x"0b",  x"3e", -- 4FA0
         x"3a",  x"cd",  x"50",  x"d2",  x"cd",  x"d2",  x"d2",  x"c3", -- 4FA8
         x"47",  x"d2",  x"fe",  x"06",  x"28",  x"0a",  x"3a",  x"58", -- 4FB0
         x"00",  x"fe",  x"12",  x"3a",  x"59",  x"00",  x"30",  x"0e", -- 4FB8
         x"06",  x"06",  x"cd",  x"41",  x"d2",  x"cd",  x"4c",  x"d0", -- 4FC0
         x"cd",  x"d2",  x"d2",  x"7b",  x"18",  x"c5",  x"f5",  x"cd", -- 4FC8
         x"0f",  x"d2",  x"fe",  x"28",  x"0e",  x"01",  x"20",  x"11", -- 4FD0
         x"0e",  x"4b",  x"f1",  x"f5",  x"fe",  x"20",  x"20",  x"04", -- 4FD8
         x"0e",  x"0a",  x"18",  x"05",  x"3e",  x"ed",  x"cd",  x"50", -- 4FE0
         x"d2",  x"79",  x"c1",  x"cd",  x"44",  x"d2",  x"18",  x"bf", -- 4FE8
         x"e1",  x"cd",  x"0f",  x"d2",  x"fe",  x"30",  x"20",  x"04", -- 4FF0
         x"3e",  x"f9",  x"18",  x"d0",  x"fe",  x"07",  x"20",  x"05", -- 4FF8
         x"cd",  x"0f",  x"d2",  x"c6",  x"10",  x"f5",  x"3e",  x"ed", -- 5000
         x"cd",  x"50",  x"d2",  x"f1",  x"18",  x"be",  x"c5",  x"cd", -- 5008
         x"0f",  x"d2",  x"20",  x"02",  x"7b",  x"3d",  x"c1",  x"c3", -- 5010
         x"44",  x"d2",  x"cd",  x"0f",  x"d2",  x"20",  x"09",  x"3e", -- 5018
         x"46",  x"80",  x"cd",  x"50",  x"d2",  x"7b",  x"18",  x"e4", -- 5020
         x"fe",  x"06",  x"28",  x"07",  x"3a",  x"58",  x"00",  x"fe", -- 5028
         x"0c",  x"30",  x"1c",  x"2b",  x"cd",  x"86",  x"00",  x"23", -- 5030
         x"fe",  x"2c",  x"28",  x"de",  x"3e",  x"05",  x"b8",  x"3a", -- 5038
         x"59",  x"00",  x"38",  x"05",  x"cd",  x"41",  x"d2",  x"18", -- 5040
         x"03",  x"cd",  x"44",  x"d2",  x"c3",  x"2d",  x"d2",  x"eb", -- 5048
         x"21",  x"d9",  x"d4",  x"78",  x"ed",  x"b1",  x"46",  x"eb", -- 5050
         x"2b",  x"cd",  x"86",  x"00",  x"23",  x"fe",  x"2c",  x"3a", -- 5058
         x"59",  x"00",  x"c2",  x"44",  x"d2",  x"78",  x"fe",  x"40", -- 5060
         x"38",  x"a4",  x"c5",  x"3e",  x"ed",  x"cd",  x"50",  x"d2", -- 5068
         x"18",  x"9d",  x"cd",  x"d2",  x"d2",  x"7b",  x"fe",  x"03", -- 5070
         x"38",  x"08",  x"3e",  x"36",  x"32",  x"80",  x"a8",  x"af", -- 5078
         x"18",  x"21",  x"11",  x"d6",  x"d4",  x"83",  x"5f",  x"1a", -- 5080
         x"18",  x"19",  x"cd",  x"0f",  x"d2",  x"4f",  x"3a",  x"59", -- 5088
         x"00",  x"3c",  x"28",  x"09",  x"cd",  x"0f",  x"d2",  x"3a", -- 5090
         x"59",  x"00",  x"3c",  x"20",  x"0b",  x"3e",  x"db",  x"cd", -- 5098
         x"50",  x"d2",  x"7b",  x"cd",  x"50",  x"d2",  x"c9",  x"4b", -- 50A0
         x"3e",  x"ed",  x"cd",  x"50",  x"d2",  x"79",  x"c3",  x"41", -- 50A8
         x"d2",  x"cd",  x"0f",  x"d2",  x"3a",  x"59",  x"00",  x"fe", -- 50B0
         x"ff",  x"f5",  x"4b",  x"cd",  x"0f",  x"d2",  x"5f",  x"f1", -- 50B8
         x"20",  x"e5",  x"3e",  x"d3",  x"cd",  x"50",  x"d2",  x"79", -- 50C0
         x"c3",  x"50",  x"d2",  x"3e",  x"cb",  x"cd",  x"50",  x"d2", -- 50C8
         x"c3",  x"b5",  x"ce",  x"cd",  x"0f",  x"d2",  x"06",  x"e3", -- 50D0
         x"fe",  x"28",  x"28",  x"11",  x"06",  x"eb",  x"fe",  x"10", -- 50D8
         x"28",  x"0b",  x"06",  x"08",  x"fe",  x"30",  x"28",  x"05", -- 50E0
         x"3e",  x"39",  x"c3",  x"e3",  x"d1",  x"c3",  x"4f",  x"d2", -- 50E8
         x"cd",  x"87",  x"d2",  x"38",  x"11",  x"fe",  x"07",  x"20", -- 50F0
         x"22",  x"2b",  x"4f",  x"cd",  x"86",  x"00",  x"23",  x"fe", -- 50F8
         x"2c",  x"79",  x"28",  x"17",  x"18",  x"0c",  x"cd",  x"0f", -- 5100
         x"d2",  x"28",  x"19",  x"3a",  x"58",  x"00",  x"fe",  x"3a", -- 5108
         x"20",  x"04",  x"06",  x"e9",  x"18",  x"d7",  x"3e",  x"41", -- 5110
         x"c3",  x"e3",  x"d1",  x"cd",  x"41",  x"d2",  x"cd",  x"d2", -- 5118
         x"d2",  x"c3",  x"47",  x"d2",  x"78",  x"06",  x"c3",  x"fe", -- 5120
         x"c2",  x"28",  x"02",  x"06",  x"cd",  x"78",  x"c3",  x"67", -- 5128
         x"cf",  x"cd",  x"87",  x"d2",  x"d2",  x"41",  x"d2",  x"cd", -- 5130
         x"d2",  x"d2",  x"20",  x"da",  x"3e",  x"c9",  x"c3",  x"50", -- 5138
         x"d2",  x"cd",  x"87",  x"d2",  x"30",  x"06",  x"78",  x"cd", -- 5140
         x"50",  x"d2",  x"18",  x"0d",  x"cb",  x"57",  x"20",  x"c6", -- 5148
         x"cb",  x"58",  x"28",  x"c2",  x"06",  x"20",  x"cd",  x"41", -- 5150
         x"d2",  x"cd",  x"0f",  x"d2",  x"20",  x"b8",  x"e5",  x"fd", -- 5158
         x"e5",  x"eb",  x"d1",  x"37",  x"ed",  x"52",  x"5d",  x"7c", -- 5160
         x"cb",  x"03",  x"ce",  x"00",  x"28",  x"0c",  x"3a",  x"80", -- 5168
         x"a8",  x"fe",  x"20",  x"20",  x"05",  x"3e",  x"36",  x"32", -- 5170
         x"80",  x"a8",  x"7d",  x"e1",  x"cd",  x"50",  x"d2",  x"c9", -- 5178
         x"cd",  x"24",  x"cb",  x"fe",  x"20",  x"30",  x"04",  x"3e", -- 5180
         x"34",  x"18",  x"58",  x"c5",  x"05",  x"20",  x"0f",  x"fe", -- 5188
         x"27",  x"20",  x"0b",  x"cd",  x"e7",  x"d1",  x"c1",  x"d8", -- 5190
         x"fe",  x"2c",  x"c0",  x"23",  x"18",  x"e2",  x"cd",  x"0f", -- 5198
         x"d2",  x"c1",  x"78",  x"fe",  x"04",  x"28",  x"13",  x"c5", -- 51A0
         x"05",  x"20",  x"01",  x"04",  x"7b",  x"cd",  x"50",  x"d2", -- 51A8
         x"7a",  x"10",  x"fa",  x"c1",  x"2b",  x"cd",  x"86",  x"00", -- 51B0
         x"18",  x"de",  x"42",  x"4b",  x"2b",  x"cd",  x"86",  x"00", -- 51B8
         x"23",  x"fe",  x"2c",  x"1e",  x"00",  x"20",  x"03",  x"cd", -- 51C0
         x"0f",  x"d2",  x"7b",  x"cd",  x"50",  x"d2",  x"0b",  x"78", -- 51C8
         x"b1",  x"20",  x"f7",  x"c9",  x"cd",  x"24",  x"cb",  x"fe", -- 51D0
         x"27",  x"20",  x"06",  x"cd",  x"e7",  x"d1",  x"fe",  x"2c", -- 51D8
         x"c0",  x"3e",  x"38",  x"32",  x"80",  x"a8",  x"c9",  x"23", -- 51E0
         x"cd",  x"86",  x"00",  x"fe",  x"20",  x"38",  x"f2",  x"23", -- 51E8
         x"fe",  x"27",  x"28",  x"05",  x"cd",  x"50",  x"d2",  x"18", -- 51F0
         x"ef",  x"cd",  x"24",  x"cb",  x"fe",  x"2c",  x"c8",  x"fe", -- 51F8
         x"3b",  x"c8",  x"fe",  x"0d",  x"c8",  x"37",  x"18",  x"d9", -- 5200
         x"cd",  x"d2",  x"d2",  x"d5",  x"fd",  x"e1",  x"c9",  x"cd", -- 5208
         x"d2",  x"d2",  x"3a",  x"54",  x"00",  x"b7",  x"28",  x"09", -- 5210
         x"32",  x"4a",  x"00",  x"3a",  x"52",  x"00",  x"32",  x"4b", -- 5218
         x"00",  x"3a",  x"55",  x"00",  x"fe",  x"28",  x"c8",  x"3a", -- 5220
         x"59",  x"00",  x"fe",  x"ff",  x"c9",  x"3a",  x"54",  x"00", -- 5228
         x"b7",  x"c8",  x"3a",  x"59",  x"00",  x"fe",  x"06",  x"37", -- 5230
         x"c0",  x"3a",  x"52",  x"00",  x"cd",  x"50",  x"d2",  x"37", -- 5238
         x"c9",  x"07",  x"07",  x"07",  x"80",  x"18",  x"09",  x"ed", -- 5240
         x"4b",  x"52",  x"00",  x"79",  x"cd",  x"50",  x"d2",  x"78", -- 5248
         x"d9",  x"4f",  x"3a",  x"3f",  x"00",  x"17",  x"17",  x"30", -- 5250
         x"08",  x"2a",  x"40",  x"00",  x"fd",  x"e5",  x"d1",  x"19", -- 5258
         x"71",  x"2a",  x"50",  x"00",  x"23",  x"22",  x"50",  x"00", -- 5260
         x"1f",  x"30",  x"18",  x"cb",  x"6f",  x"28",  x"05",  x"cd", -- 5268
         x"fb",  x"d6",  x"18",  x"0f",  x"3e",  x"8f",  x"2a",  x"48", -- 5270
         x"00",  x"bd",  x"28",  x"07",  x"79",  x"cd",  x"b7",  x"cb", -- 5278
         x"22",  x"48",  x"00",  x"d9",  x"fd",  x"23",  x"c9",  x"c5", -- 5280
         x"e5",  x"cd",  x"24",  x"cb",  x"cd",  x"89",  x"d6",  x"38", -- 5288
         x"3d",  x"57",  x"1e",  x"20",  x"23",  x"cd",  x"86",  x"00", -- 5290
         x"cd",  x"75",  x"d6",  x"38",  x"0a",  x"5f",  x"23",  x"cd", -- 5298
         x"86",  x"00",  x"cd",  x"75",  x"d6",  x"30",  x"27",  x"cd", -- 52A0
         x"24",  x"cb",  x"fe",  x"2c",  x"20",  x"01",  x"23",  x"e5", -- 52A8
         x"21",  x"f2",  x"d4",  x"01",  x"10",  x"00",  x"7b",  x"ed", -- 52B0
         x"b9",  x"20",  x"12",  x"7a",  x"be",  x"28",  x"04",  x"79", -- 52B8
         x"b7",  x"20",  x"f3",  x"cb",  x"39",  x"30",  x"06",  x"79", -- 52C0
         x"e1",  x"d1",  x"c1",  x"3f",  x"c9",  x"e1",  x"e1",  x"c1", -- 52C8
         x"37",  x"c9",  x"c5",  x"af",  x"d9",  x"06",  x"08",  x"21", -- 52D0
         x"51",  x"00",  x"23",  x"77",  x"10",  x"fc",  x"35",  x"d9", -- 52D8
         x"3e",  x"2b",  x"32",  x"57",  x"00",  x"2b",  x"23",  x"cd", -- 52E0
         x"24",  x"cb",  x"fe",  x"3b",  x"28",  x"3c",  x"fe",  x"20", -- 52E8
         x"38",  x"38",  x"32",  x"56",  x"00",  x"fe",  x"27",  x"ca", -- 52F0
         x"84",  x"d3",  x"fe",  x"2c",  x"28",  x"2b",  x"fe",  x"28", -- 52F8
         x"28",  x"32",  x"fe",  x"29",  x"28",  x"e0",  x"fe",  x"2d", -- 5300
         x"28",  x"2f",  x"fe",  x"2b",  x"28",  x"2b",  x"fe",  x"2a", -- 5308
         x"28",  x"27",  x"fe",  x"2f",  x"28",  x"23",  x"fe",  x"25", -- 5310
         x"28",  x"1f",  x"fe",  x"24",  x"28",  x"04",  x"fe",  x"23", -- 5318
         x"20",  x"1c",  x"ed",  x"4b",  x"4c",  x"00",  x"c3",  x"a6", -- 5320
         x"d3",  x"23",  x"ed",  x"5b",  x"52",  x"00",  x"c1",  x"3a", -- 5328
         x"56",  x"00",  x"b7",  x"c9",  x"32",  x"55",  x"00",  x"18", -- 5330
         x"ad",  x"32",  x"57",  x"00",  x"18",  x"a8",  x"cd",  x"89", -- 5338
         x"d6",  x"d2",  x"3d",  x"d4",  x"e5",  x"0e",  x"0a",  x"cd", -- 5340
         x"18",  x"d6",  x"38",  x"08",  x"e1",  x"23",  x"e5",  x"3e", -- 5348
         x"35",  x"32",  x"80",  x"a8",  x"0e",  x"10",  x"cd",  x"18", -- 5350
         x"d6",  x"38",  x"fb",  x"e1",  x"fe",  x"11",  x"28",  x"02", -- 5358
         x"0e",  x"0a",  x"e5",  x"21",  x"00",  x"00",  x"e3",  x"cd", -- 5360
         x"18",  x"d6",  x"e3",  x"38",  x"0b",  x"fe",  x"11",  x"28", -- 5368
         x"03",  x"e3",  x"2b",  x"e3",  x"d5",  x"c1",  x"18",  x"5f", -- 5370
         x"5f",  x"af",  x"57",  x"19",  x"eb",  x"6f",  x"41",  x"19", -- 5378
         x"10",  x"fd",  x"18",  x"e2",  x"01",  x"00",  x"00",  x"3a", -- 5380
         x"58",  x"00",  x"fe",  x"2d",  x"ca",  x"e6",  x"d2",  x"23", -- 5388
         x"cd",  x"86",  x"00",  x"fe",  x"27",  x"28",  x"0f",  x"fe", -- 5390
         x"20",  x"38",  x"04",  x"41",  x"4f",  x"18",  x"f0",  x"3e", -- 5398
         x"38",  x"32",  x"80",  x"a8",  x"18",  x"01",  x"23",  x"e5", -- 53A0
         x"18",  x"2d",  x"f1",  x"1b",  x"1b",  x"eb",  x"cd",  x"2d", -- 53A8
         x"d6",  x"d5",  x"2b",  x"cd",  x"86",  x"00",  x"3d",  x"20", -- 53B0
         x"05",  x"3e",  x"32",  x"32",  x"80",  x"a8",  x"2b",  x"cd", -- 53B8
         x"86",  x"00",  x"47",  x"2b",  x"cd",  x"86",  x"00",  x"4f", -- 53C0
         x"30",  x"0d",  x"e1",  x"cd",  x"39",  x"cb",  x"d5",  x"3e", -- 53C8
         x"33",  x"32",  x"80",  x"a8",  x"01",  x"00",  x"00",  x"21", -- 53D0
         x"57",  x"00",  x"7e",  x"36",  x"00",  x"2a",  x"52",  x"00", -- 53D8
         x"fe",  x"2b",  x"28",  x"1c",  x"fe",  x"2d",  x"28",  x"1b", -- 53E0
         x"fe",  x"2a",  x"28",  x"1b",  x"fe",  x"2f",  x"28",  x"32", -- 53E8
         x"fe",  x"25",  x"28",  x"33",  x"3e",  x"42",  x"32",  x"80", -- 53F0
         x"a8",  x"22",  x"52",  x"00",  x"e1",  x"c3",  x"e7",  x"d2", -- 53F8
         x"09",  x"18",  x"f6",  x"ed",  x"42",  x"18",  x"f2",  x"eb", -- 5400
         x"21",  x"00",  x"00",  x"3e",  x"10",  x"cb",  x"1a",  x"cb", -- 5408
         x"1b",  x"30",  x"01",  x"09",  x"cb",  x"1c",  x"cb",  x"1d", -- 5410
         x"cb",  x"1a",  x"cb",  x"1b",  x"3d",  x"20",  x"f2",  x"eb", -- 5418
         x"18",  x"d7",  x"cd",  x"2c",  x"d4",  x"18",  x"f8",  x"cd", -- 5420
         x"2c",  x"d4",  x"18",  x"cd",  x"11",  x"ff",  x"ff",  x"78", -- 5428
         x"b1",  x"3e",  x"43",  x"ca",  x"e3",  x"d1",  x"13",  x"ed", -- 5430
         x"42",  x"30",  x"fb",  x"09",  x"c9",  x"f5",  x"23",  x"cd", -- 5438
         x"86",  x"00",  x"eb",  x"cd",  x"75",  x"d6",  x"30",  x"24", -- 5440
         x"f1",  x"fe",  x"4d",  x"20",  x"10",  x"cd",  x"8c",  x"00", -- 5448
         x"fe",  x"30",  x"d2",  x"ac",  x"d3",  x"3e",  x"28",  x"32", -- 5450
         x"55",  x"00",  x"eb",  x"18",  x"75",  x"21",  x"03",  x"d5", -- 5458
         x"01",  x"09",  x"00",  x"ed",  x"b1",  x"c2",  x"ac",  x"d3", -- 5460
         x"cb",  x"21",  x"18",  x"29",  x"13",  x"21",  x"1a",  x"d5", -- 5468
         x"01",  x"16",  x"00",  x"ed",  x"a9",  x"28",  x"07",  x"ed", -- 5470
         x"a9",  x"e2",  x"aa",  x"d3",  x"18",  x"f5",  x"47",  x"cd", -- 5478
         x"8c",  x"00",  x"cd",  x"75",  x"d6",  x"d2",  x"aa",  x"d3", -- 5480
         x"f1",  x"be",  x"28",  x"06",  x"f5",  x"78",  x"06",  x"00", -- 5488
         x"18",  x"e5",  x"80",  x"d6",  x"19",  x"d6",  x"41",  x"06", -- 5490
         x"00",  x"eb",  x"32",  x"58",  x"00",  x"fe",  x"3a",  x"20", -- 5498
         x"14",  x"3a",  x"55",  x"00",  x"b7",  x"3e",  x"20",  x"28", -- 54A0
         x"06",  x"af",  x"32",  x"55",  x"00",  x"3e",  x"06",  x"32", -- 54A8
         x"59",  x"00",  x"c3",  x"e7",  x"d2",  x"e5",  x"21",  x"1b", -- 54B0
         x"d5",  x"09",  x"7e",  x"e1",  x"b7",  x"f2",  x"af",  x"d4", -- 54B8
         x"f5",  x"f6",  x"0d",  x"32",  x"54",  x"00",  x"f1",  x"e6", -- 54C0
         x"0f",  x"fe",  x"0d",  x"28",  x"05",  x"f6",  x"40",  x"eb", -- 54C8
         x"18",  x"8b",  x"3e",  x"3a",  x"18",  x"c4",  x"46",  x"56", -- 54D0
         x"5e",  x"05",  x"0b",  x"04",  x"03",  x"80",  x"09",  x"88", -- 54D8
         x"4a",  x"98",  x"42",  x"4e",  x"5a",  x"5a",  x"20",  x"4e", -- 54E0
         x"43",  x"43",  x"20",  x"50",  x"4f",  x"50",  x"45",  x"50", -- 54E8
         x"20",  x"4d",  x"20",  x"00",  x"09",  x"6f",  x"fd",  x"0c", -- 54F0
         x"58",  x"18",  x"27",  x"1a",  x"08",  x"1d",  x"41",  x"10", -- 54F8
         x"3f",  x"54",  x"34",  x"49",  x"52",  x"42",  x"43",  x"44", -- 5500
         x"45",  x"48",  x"4c",  x"41",  x"46",  x"53",  x"50",  x"49", -- 5508
         x"58",  x"49",  x"59",  x"48",  x"58",  x"48",  x"59",  x"4c", -- 5510
         x"58",  x"4c",  x"59",  x"07",  x"00",  x"05",  x"10",  x"04", -- 5518
         x"20",  x"03",  x"30",  x"02",  x"30",  x"01",  x"dd",  x"00", -- 5520
         x"fd",  x"4f",  x"d8",  x"47",  x"f8",  x"ff",  x"dc",  x"ff", -- 5528
         x"fc",  x"40",  x"b8",  x"40",  x"c2",  x"45",  x"38",  x"28", -- 5530
         x"18",  x"88",  x"80",  x"c4",  x"18",  x"05",  x"f4",  x"fc", -- 5538
         x"40",  x"00",  x"02",  x"70",  x"a0",  x"a9",  x"b9",  x"47", -- 5540
         x"aa",  x"98",  x"a1",  x"04",  x"ab",  x"a2",  x"00",  x"10", -- 5548
         x"30",  x"20",  x"b0",  x"08",  x"68",  x"18",  x"20",  x"28", -- 5550
         x"08",  x"10",  x"77",  x"80",  x"c0",  x"c0",  x"01",  x"b2", -- 5558
         x"c1",  x"00",  x"38",  x"30",  x"ba",  x"4e",  x"da",  x"10", -- 5560
         x"b1",  x"41",  x"46",  x"bb",  x"c8",  x"ac",  x"a3",  x"b4", -- 5568
         x"bc",  x"c5",  x"a4",  x"a8",  x"00",  x"00",  x"03",  x"90", -- 5570
         x"01",  x"03",  x"04",  x"04",  x"b3",  x"00",  x"72",  x"71", -- 5578
         x"43",  x"34",  x"76",  x"2a",  x"a3",  x"43",  x"33",  x"4c", -- 5580
         x"74",  x"04",  x"4a",  x"73",  x"54",  x"13",  x"33",  x"71", -- 5588
         x"42",  x"2d",  x"a3",  x"44",  x"c3",  x"e3",  x"f5",  x"83", -- 5590
         x"34",  x"93",  x"34",  x"c3",  x"d3",  x"29",  x"08",  x"03", -- 5598
         x"58",  x"04",  x"73",  x"83",  x"68",  x"53",  x"18",  x"78", -- 55A0
         x"73",  x"03",  x"51",  x"6b",  x"21",  x"63",  x"c3",  x"63", -- 55A8
         x"0f",  x"48",  x"78",  x"93",  x"d3",  x"43",  x"6c",  x"b3", -- 55B0
         x"27",  x"a3",  x"d3",  x"13",  x"83",  x"83",  x"c3",  x"93", -- 55B8
         x"23",  x"d3",  x"14",  x"4e",  x"18",  x"6d",  x"24",  x"6d", -- 55C0
         x"3d",  x"7d",  x"2d",  x"a3",  x"70",  x"a3",  x"d3",  x"a2", -- 55C8
         x"e2",  x"18",  x"16",  x"20",  x"8c",  x"7d",  x"58",  x"26", -- 55D0
         x"40",  x"4d",  x"61",  x"2e",  x"89",  x"63",  x"64",  x"8a", -- 55D8
         x"57",  x"98",  x"67",  x"72",  x"78",  x"94",  x"9a",  x"82", -- 55E0
         x"90",  x"0a",  x"8b",  x"1b",  x"75",  x"a4",  x"34",  x"46", -- 55E8
         x"24",  x"1f",  x"49",  x"65",  x"70",  x"53",  x"da",  x"4d", -- 55F0
         x"3f",  x"00",  x"01",  x"02",  x"03",  x"04",  x"05",  x"07", -- 55F8
         x"0a",  x"43",  x"0b",  x"0f",  x"3d",  x"44",  x"12",  x"15", -- 5600
         x"45",  x"23",  x"30",  x"33",  x"46",  x"37",  x"3a",  x"3b", -- 5608
         x"42",  x"47",  x"48",  x"49",  x"4a",  x"4b",  x"4c",  x"4e", -- 5610
         x"cd",  x"86",  x"00",  x"cd",  x"89",  x"d6",  x"23",  x"fe", -- 5618
         x"3a",  x"30",  x"02",  x"d6",  x"30",  x"fe",  x"41",  x"38", -- 5620
         x"02",  x"d6",  x"37",  x"b9",  x"c9",  x"e5",  x"2a",  x"44", -- 5628
         x"00",  x"e5",  x"ed",  x"5b",  x"46",  x"00",  x"1b",  x"b7", -- 5630
         x"ed",  x"52",  x"44",  x"4d",  x"e1",  x"d1",  x"cd",  x"8c", -- 5638
         x"00",  x"cd",  x"89",  x"d6",  x"cd",  x"78",  x"00",  x"37", -- 5640
         x"e0",  x"cd",  x"31",  x"cb",  x"38",  x"f0",  x"c9",  x"21", -- 5648
         x"5a",  x"cc",  x"11",  x"23",  x"00",  x"01",  x"06",  x"00", -- 5650
         x"ed",  x"b0",  x"21",  x"23",  x"00",  x"cd",  x"2d",  x"d6", -- 5658
         x"d8",  x"2b",  x"cd",  x"86",  x"00",  x"3d",  x"37",  x"c8", -- 5660
         x"2b",  x"cd",  x"86",  x"00",  x"f5",  x"2b",  x"cd",  x"86", -- 5668
         x"00",  x"e1",  x"6f",  x"a7",  x"c9",  x"cd",  x"89",  x"d6", -- 5670
         x"d0",  x"fe",  x"30",  x"38",  x"04",  x"fe",  x"3a",  x"3f", -- 5678
         x"d0",  x"fe",  x"2e",  x"c8",  x"fe",  x"5f",  x"c8",  x"37", -- 5680
         x"c9",  x"fe",  x"41",  x"d8",  x"fe",  x"5b",  x"3f",  x"d0", -- 5688
         x"fe",  x"61",  x"d8",  x"fe",  x"7b",  x"3f",  x"d8",  x"e6", -- 5690
         x"df",  x"c9",  x"c5",  x"06",  x"01",  x"fe",  x"20",  x"30", -- 5698
         x"21",  x"fe",  x"0c",  x"28",  x"09",  x"fe",  x"0d",  x"20", -- 56A0
         x"09",  x"cd",  x"55",  x"c5",  x"3e",  x"0a",  x"1e",  x"ff", -- 56A8
         x"18",  x"10",  x"fe",  x"09",  x"20",  x"16",  x"3e",  x"08", -- 56B0
         x"93",  x"e6",  x"07",  x"20",  x"02",  x"3e",  x"08",  x"47", -- 56B8
         x"3e",  x"20",  x"cd",  x"55",  x"c5",  x"1c",  x"7b",  x"ba", -- 56C0
         x"28",  x"02",  x"10",  x"f4",  x"cd",  x"d1",  x"c7",  x"c1", -- 56C8
         x"c9",  x"cd",  x"03",  x"f0",  x"20",  x"11",  x"d1",  x"c8", -- 56D0
         x"cd",  x"8b",  x"c8",  x"30",  x"03",  x"e1",  x"e1",  x"c9", -- 56D8
         x"cd",  x"d5",  x"c8",  x"3e",  x"02",  x"32",  x"10",  x"b7", -- 56E0
         x"2a",  x"50",  x"00",  x"22",  x"13",  x"b7",  x"cd",  x"4f", -- 56E8
         x"d6",  x"d8",  x"3e",  x"03",  x"32",  x"10",  x"b7",  x"22", -- 56F0
         x"15",  x"b7",  x"c9",  x"c5",  x"21",  x"3e",  x"00",  x"cb", -- 56F8
         x"5e",  x"28",  x"4e",  x"cb",  x"9e",  x"21",  x"00",  x"b7", -- 5700
         x"dd",  x"75",  x"05",  x"dd",  x"74",  x"06",  x"fd",  x"e5", -- 5708
         x"d1",  x"2a",  x"13",  x"b7",  x"19",  x"ed",  x"53",  x"11", -- 5710
         x"b7",  x"22",  x"13",  x"b7",  x"eb",  x"cd",  x"03",  x"f0", -- 5718
         x"1b",  x"3a",  x"10",  x"b7",  x"fe",  x"03",  x"38",  x"07", -- 5720
         x"2a",  x"15",  x"b7",  x"cd",  x"03",  x"f0",  x"1a",  x"cd", -- 5728
         x"50",  x"c5",  x"21",  x"00",  x"b7",  x"cd",  x"03",  x"f0", -- 5730
         x"08",  x"08",  x"21",  x"80",  x"b7",  x"af",  x"2d",  x"77", -- 5738
         x"20",  x"fc",  x"08",  x"dd",  x"7e",  x"02",  x"cd",  x"03", -- 5740
         x"f0",  x"1c",  x"cd",  x"03",  x"f0",  x"23",  x"08",  x"08", -- 5748
         x"00",  x"21",  x"00",  x"b7",  x"08",  x"fe",  x"80",  x"20", -- 5750
         x"09",  x"01",  x"a0",  x"00",  x"cd",  x"03",  x"f0",  x"01", -- 5758
         x"18",  x"d8",  x"6f",  x"3c",  x"08",  x"c1",  x"71",  x"c9", -- 5760
         x"dd",  x"dd",  x"44",  x"49",  x"52",  x"1f",  x"cd",  x"21", -- 5768
         x"f0",  x"08",  x"c9",  x"dd",  x"dd",  x"43",  x"44",  x"1f", -- 5770
         x"cd",  x"21",  x"f0",  x"09",  x"c9",  x"dd",  x"dd",  x"52", -- 5778
         x"45",  x"4e",  x"1f",  x"cd",  x"21",  x"f0",  x"0b",  x"c9", -- 5780
         x"dd",  x"dd",  x"45",  x"52",  x"41",  x"1f",  x"cd",  x"21", -- 5788
         x"f0",  x"0a",  x"c9",  x"dd",  x"dd",  x"44",  x"45",  x"56", -- 5790
         x"49",  x"43",  x"45",  x"01",  x"a7",  x"28",  x"0e",  x"7d", -- 5798
         x"fe",  x"08",  x"30",  x"04",  x"cd",  x"af",  x"d7",  x"d0", -- 57A0
         x"cd",  x"03",  x"f0",  x"19",  x"c9",  x"3e",  x"ff",  x"cd", -- 57A8
         x"03",  x"f0",  x"49",  x"c9",  x"7f",  x"7f",  x"53",  x"45", -- 57B0
         x"54",  x"52",  x"4f",  x"1f",  x"21",  x"52",  x"d9",  x"e5", -- 57B8
         x"cd",  x"1c",  x"d8",  x"cd",  x"5d",  x"d8",  x"3e",  x"25", -- 57C0
         x"18",  x"14",  x"7f",  x"7f",  x"53",  x"45",  x"54",  x"57", -- 57C8
         x"52",  x"1f",  x"21",  x"52",  x"d9",  x"e5",  x"cd",  x"1c", -- 57D0
         x"d8",  x"cd",  x"5d",  x"d8",  x"3e",  x"31",  x"d8",  x"01", -- 57D8
         x"f3",  x"80",  x"ed",  x"79",  x"c5",  x"3e",  x"01",  x"cd", -- 57E0
         x"03",  x"f0",  x"14",  x"c1",  x"ed",  x"78",  x"a7",  x"cb", -- 57E8
         x"47",  x"20",  x"f1",  x"cb",  x"7f",  x"c8",  x"01",  x"f1", -- 57F0
         x"83",  x"ed",  x"78",  x"fe",  x"20",  x"30",  x"0f",  x"01", -- 57F8
         x"f3",  x"81",  x"ed",  x"78",  x"cd",  x"03",  x"f0",  x"1c", -- 5800
         x"cd",  x"03",  x"f0",  x"19",  x"37",  x"c9",  x"06",  x"00", -- 5808
         x"ed",  x"78",  x"04",  x"a7",  x"28",  x"f6",  x"cd",  x"03", -- 5810
         x"f0",  x"24",  x"18",  x"f4",  x"01",  x"80",  x"fc",  x"ed", -- 5818
         x"78",  x"fe",  x"a7",  x"28",  x"14",  x"cd",  x"03",  x"f0", -- 5820
         x"23",  x"4b",  x"65",  x"69",  x"6e",  x"20",  x"44",  x"30", -- 5828
         x"30",  x"34",  x"21",  x"07",  x"0d",  x"0a",  x"00",  x"e1", -- 5830
         x"c9",  x"01",  x"f3",  x"b3",  x"ed",  x"78",  x"fe",  x"05", -- 5838
         x"c8",  x"cd",  x"03",  x"f0",  x"23",  x"43",  x"41",  x"4f", -- 5840
         x"53",  x"2d",  x"44",  x"69",  x"73",  x"6b",  x"20",  x"73", -- 5848
         x"74",  x"61",  x"72",  x"74",  x"65",  x"6e",  x"21",  x"07", -- 5850
         x"0d",  x"0a",  x"00",  x"e1",  x"c9",  x"eb",  x"7e",  x"e6", -- 5858
         x"df",  x"20",  x"14",  x"21",  x"06",  x"00",  x"cd",  x"03", -- 5860
         x"f0",  x"23",  x"4e",  x"61",  x"6d",  x"65",  x"20",  x"3a", -- 5868
         x"00",  x"cd",  x"03",  x"f0",  x"17",  x"d8",  x"19",  x"1e", -- 5870
         x"0c",  x"01",  x"f3",  x"82",  x"7e",  x"ed",  x"79",  x"e6", -- 5878
         x"df",  x"28",  x"01",  x"23",  x"04",  x"1d",  x"20",  x"f4", -- 5880
         x"eb",  x"13",  x"c9",  x"7f",  x"7f",  x"54",  x"49",  x"4d", -- 5888
         x"45",  x"01",  x"21",  x"52",  x"d9",  x"e5",  x"cd",  x"1c", -- 5890
         x"d8",  x"01",  x"f1",  x"83",  x"ed",  x"78",  x"fe",  x"30", -- 5898
         x"30",  x"14",  x"cd",  x"03",  x"f0",  x"23",  x"4b",  x"65", -- 58A0
         x"69",  x"6e",  x"20",  x"44",  x"45",  x"50",  x"20",  x"33", -- 58A8
         x"21",  x"07",  x"0d",  x"0a",  x"00",  x"c9",  x"3e",  x"19", -- 58B0
         x"cd",  x"03",  x"f0",  x"24",  x"1e",  x"02",  x"01",  x"f1", -- 58B8
         x"86",  x"ed",  x"78",  x"cd",  x"03",  x"f0",  x"1c",  x"3e", -- 58C0
         x"2e",  x"cd",  x"03",  x"f0",  x"24",  x"05",  x"1d",  x"20", -- 58C8
         x"f0",  x"ed",  x"78",  x"fe",  x"78",  x"3e",  x"19",  x"ce", -- 58D0
         x"00",  x"27",  x"cd",  x"03",  x"f0",  x"1c",  x"ed",  x"78", -- 58D8
         x"cd",  x"03",  x"f0",  x"1c",  x"cd",  x"03",  x"f0",  x"23", -- 58E0
         x"20",  x"00",  x"1e",  x"02",  x"01",  x"f1",  x"87",  x"ed", -- 58E8
         x"78",  x"cd",  x"03",  x"f0",  x"1c",  x"3e",  x"3a",  x"cd", -- 58F0
         x"03",  x"f0",  x"24",  x"04",  x"1d",  x"20",  x"f0",  x"ed", -- 58F8
         x"78",  x"cd",  x"03",  x"f0",  x"1c",  x"3a",  x"81",  x"b7", -- 5900
         x"a7",  x"28",  x"06",  x"cd",  x"03",  x"f0",  x"2a",  x"30", -- 5908
         x"a5",  x"cd",  x"03",  x"f0",  x"2c",  x"c9",  x"7f",  x"7f", -- 5910
         x"50",  x"52",  x"49",  x"4e",  x"54",  x"1f",  x"21",  x"52", -- 5918
         x"d9",  x"e5",  x"1a",  x"a7",  x"c8",  x"fe",  x"20",  x"28", -- 5920
         x"15",  x"fe",  x"2c",  x"28",  x"14",  x"fe",  x"27",  x"28", -- 5928
         x"14",  x"cd",  x"03",  x"f0",  x"18",  x"da",  x"19",  x"00", -- 5930
         x"3a",  x"97",  x"b7",  x"cd",  x"e9",  x"b7",  x"13",  x"18", -- 5938
         x"e1",  x"13",  x"1a",  x"18",  x"f6",  x"13",  x"1a",  x"a7", -- 5940
         x"c8",  x"fe",  x"27",  x"28",  x"f1",  x"cd",  x"e9",  x"b7", -- 5948
         x"18",  x"f3",  x"ed",  x"5b",  x"7f",  x"b7",  x"3e",  x"02", -- 5950
         x"6f",  x"1e",  x"26",  x"c3",  x"09",  x"f0",  x"ff",  x"ff", -- 5958
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5960
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5968
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5970
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5978
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5980
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5988
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5990
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5998
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 59A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 59A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 59B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 59B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 59C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 59C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 59D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 59D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 59E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 59E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 59F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 59F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5A98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5AA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5AA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5AB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5AB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5AC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5AC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5AD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5AD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5AE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5AE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5AF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5AF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5B98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5BA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5BA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5BB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5BB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5BC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5BC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5BD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5BD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5BE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5BE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5BF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5BF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5C98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5CA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5CA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5CB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5CB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5CC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5CC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5CD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5CD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5CE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5CE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5CF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5CF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5D98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5DA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5DA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5DB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5DB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5DC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5DC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5DD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5DD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5DE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5DE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5DF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5DF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5E98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5EA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5EA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5EB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5EB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5EC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5EC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5ED0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5ED8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5EE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5EE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5EF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5EF8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F00
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F08
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F10
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F18
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F20
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F28
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F30
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F38
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F40
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F48
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F50
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F58
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F60
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F68
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F70
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F78
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F80
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F88
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F90
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5F98
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5FA0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5FA8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5FB0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5FB8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5FC0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5FC8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5FD0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5FD8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5FE0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5FE8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5FF0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 5FF8
         x"18",  x"0b",  x"c3",  x"8c",  x"c0",  x"7f",  x"7f",  x"42", -- 6000
         x"41",  x"53",  x"49",  x"43",  x"00",  x"21",  x"bd",  x"c0", -- 6008
         x"11",  x"00",  x"03",  x"01",  x"67",  x"00",  x"ed",  x"b0", -- 6010
         x"eb",  x"f9",  x"cd",  x"69",  x"c6",  x"32",  x"ab",  x"03", -- 6018
         x"32",  x"00",  x"04",  x"21",  x"92",  x"c0",  x"cd",  x"c9", -- 6020
         x"d1",  x"21",  x"ae",  x"c0",  x"cd",  x"c9",  x"d1",  x"cd", -- 6028
         x"ae",  x"c5",  x"21",  x"62",  x"03",  x"cd",  x"86",  x"c9", -- 6030
         x"7a",  x"d6",  x"06",  x"21",  x"00",  x"03",  x"2b",  x"30", -- 6038
         x"03",  x"11",  x"ff",  x"bf",  x"23",  x"cd",  x"89",  x"c6", -- 6040
         x"28",  x"09",  x"7e",  x"47",  x"2f",  x"77",  x"be",  x"70", -- 6048
         x"28",  x"f2",  x"2b",  x"11",  x"00",  x"ff",  x"22",  x"b0", -- 6050
         x"03",  x"19",  x"22",  x"56",  x"03",  x"cd",  x"41",  x"c6", -- 6058
         x"2a",  x"56",  x"03",  x"11",  x"ef",  x"fb",  x"19",  x"cd", -- 6060
         x"29",  x"d8",  x"21",  x"a0",  x"c0",  x"cd",  x"c9",  x"d1", -- 6068
         x"2a",  x"04",  x"e0",  x"7e",  x"fe",  x"78",  x"20",  x"01", -- 6070
         x"3e",  x"af",  x"32",  x"fc",  x"03",  x"31",  x"67",  x"03", -- 6078
         x"18",  x"0a",  x"7f",  x"7f",  x"52",  x"45",  x"42",  x"41", -- 6080
         x"53",  x"49",  x"43",  x"00",  x"cd",  x"69",  x"c6",  x"c3", -- 6088
         x"88",  x"c3",  x"0c",  x"0a",  x"0d",  x"48",  x"43",  x"2d", -- 6090
         x"42",  x"41",  x"53",  x"49",  x"43",  x"0a",  x"0d",  x"00", -- 6098
         x"20",  x"42",  x"59",  x"54",  x"45",  x"53",  x"20",  x"46", -- 60A0
         x"52",  x"45",  x"45",  x"0a",  x"0d",  x"00",  x"4d",  x"45", -- 60A8
         x"4d",  x"4f",  x"52",  x"59",  x"20",  x"45",  x"4e",  x"44", -- 60B0
         x"20",  x"3f",  x"20",  x"3a",  x"00",  x"c3",  x"89",  x"c0", -- 60B8
         x"c3",  x"67",  x"c9",  x"00",  x"00",  x"00",  x"00",  x"00", -- 60C0
         x"d6",  x"00",  x"6f",  x"7c",  x"de",  x"00",  x"67",  x"78", -- 60C8
         x"de",  x"00",  x"47",  x"3e",  x"00",  x"c9",  x"00",  x"00", -- 60D0
         x"00",  x"35",  x"4a",  x"ca",  x"99",  x"39",  x"1c",  x"76", -- 60D8
         x"98",  x"22",  x"95",  x"b3",  x"98",  x"0a",  x"dd",  x"47", -- 60E0
         x"98",  x"53",  x"d1",  x"99",  x"99",  x"0a",  x"1a",  x"9f", -- 60E8
         x"98",  x"65",  x"bc",  x"cd",  x"98",  x"d6",  x"77",  x"3e", -- 60F0
         x"98",  x"52",  x"c7",  x"4f",  x"80",  x"0b",  x"ff",  x"1b", -- 60F8
         x"00",  x"0a",  x"00",  x"0a",  x"00",  x"00",  x"00",  x"c3", -- 6100
         x"ae",  x"c5",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 6108
         x"00",  x"00",  x"00",  x"65",  x"04",  x"fe",  x"ff",  x"00", -- 6110
         x"00",  x"c9",  x"00",  x"00",  x"01",  x"04",  x"00",  x"00", -- 6118
         x"00",  x"c5",  x"4e",  x"44",  x"c6",  x"4f",  x"52",  x"ce", -- 6120
         x"45",  x"58",  x"54",  x"c4",  x"41",  x"54",  x"41",  x"c9", -- 6128
         x"4e",  x"50",  x"55",  x"54",  x"c4",  x"49",  x"4d",  x"d2", -- 6130
         x"45",  x"41",  x"44",  x"cc",  x"45",  x"54",  x"c7",  x"4f", -- 6138
         x"54",  x"4f",  x"d2",  x"55",  x"4e",  x"c9",  x"46",  x"d2", -- 6140
         x"45",  x"53",  x"54",  x"4f",  x"52",  x"45",  x"c7",  x"4f", -- 6148
         x"53",  x"55",  x"42",  x"d2",  x"45",  x"54",  x"55",  x"52", -- 6150
         x"4e",  x"d2",  x"45",  x"4d",  x"d3",  x"54",  x"4f",  x"50", -- 6158
         x"cf",  x"55",  x"54",  x"cf",  x"4e",  x"ce",  x"55",  x"4c", -- 6160
         x"4c",  x"d7",  x"41",  x"49",  x"54",  x"c4",  x"45",  x"46", -- 6168
         x"d0",  x"4f",  x"4b",  x"45",  x"c4",  x"4f",  x"4b",  x"45", -- 6170
         x"c1",  x"55",  x"54",  x"4f",  x"cc",  x"49",  x"4e",  x"45", -- 6178
         x"53",  x"c3",  x"4c",  x"53",  x"d7",  x"49",  x"44",  x"54", -- 6180
         x"48",  x"c2",  x"59",  x"45",  x"a1",  x"c3",  x"41",  x"4c", -- 6188
         x"4c",  x"d0",  x"52",  x"49",  x"4e",  x"54",  x"c3",  x"4f", -- 6190
         x"4e",  x"54",  x"cc",  x"49",  x"53",  x"54",  x"c3",  x"4c", -- 6198
         x"45",  x"41",  x"52",  x"c3",  x"4c",  x"4f",  x"41",  x"44", -- 61A0
         x"c3",  x"53",  x"41",  x"56",  x"45",  x"ce",  x"45",  x"57", -- 61A8
         x"d4",  x"41",  x"42",  x"28",  x"d4",  x"4f",  x"c6",  x"4e", -- 61B0
         x"d3",  x"50",  x"43",  x"28",  x"d4",  x"48",  x"45",  x"4e", -- 61B8
         x"ce",  x"4f",  x"54",  x"d3",  x"54",  x"45",  x"50",  x"ab", -- 61C0
         x"ad",  x"aa",  x"af",  x"de",  x"c1",  x"4e",  x"44",  x"cf", -- 61C8
         x"52",  x"be",  x"bd",  x"bc",  x"d3",  x"47",  x"4e",  x"c9", -- 61D0
         x"4e",  x"54",  x"c1",  x"42",  x"53",  x"d5",  x"53",  x"52", -- 61D8
         x"c6",  x"52",  x"45",  x"c9",  x"4e",  x"50",  x"d0",  x"4f", -- 61E0
         x"53",  x"d3",  x"51",  x"52",  x"d2",  x"4e",  x"44",  x"cc", -- 61E8
         x"4e",  x"c5",  x"58",  x"50",  x"c3",  x"4f",  x"53",  x"d3", -- 61F0
         x"49",  x"4e",  x"d4",  x"41",  x"4e",  x"c1",  x"54",  x"4e", -- 61F8
         x"d0",  x"45",  x"45",  x"4b",  x"c4",  x"45",  x"45",  x"4b", -- 6200
         x"d0",  x"49",  x"cc",  x"45",  x"4e",  x"d3",  x"54",  x"52", -- 6208
         x"24",  x"d6",  x"41",  x"4c",  x"c1",  x"53",  x"43",  x"c3", -- 6210
         x"48",  x"52",  x"24",  x"cc",  x"45",  x"46",  x"54",  x"24", -- 6218
         x"d2",  x"49",  x"47",  x"48",  x"54",  x"24",  x"cd",  x"49", -- 6220
         x"44",  x"24",  x"cc",  x"4f",  x"41",  x"44",  x"d4",  x"52", -- 6228
         x"4f",  x"4e",  x"d4",  x"52",  x"4f",  x"46",  x"46",  x"c5", -- 6230
         x"44",  x"49",  x"54",  x"c5",  x"4c",  x"53",  x"45",  x"80", -- 6238
         x"1a",  x"c9",  x"de",  x"c7",  x"dc",  x"cc",  x"48",  x"ca", -- 6240
         x"ec",  x"cb",  x"01",  x"cf",  x"1f",  x"cc",  x"5d",  x"ca", -- 6248
         x"07",  x"ca",  x"eb",  x"c9",  x"cf",  x"ca",  x"df",  x"c8", -- 6250
         x"f6",  x"c9",  x"25",  x"ca",  x"4a",  x"ca",  x"18",  x"c9", -- 6258
         x"ec",  x"d3",  x"b3",  x"ca",  x"c0",  x"cb",  x"f7",  x"d3", -- 6260
         x"c4",  x"d0",  x"37",  x"d4",  x"4e",  x"d4",  x"fa",  x"c5", -- 6268
         x"ea",  x"c6",  x"d0",  x"dd",  x"b9",  x"cb",  x"f4",  x"df", -- 6270
         x"4a",  x"ca",  x"38",  x"db",  x"fa",  x"ca",  x"48",  x"c9", -- 6278
         x"f2",  x"c6",  x"aa",  x"c9",  x"43",  x"dc",  x"41",  x"dd", -- 6280
         x"40",  x"c6",  x"2d",  x"c6",  x"b7",  x"c7",  x"b8",  x"c7", -- 6288
         x"e7",  x"c3",  x"4a",  x"ca",  x"a6",  x"d6",  x"70",  x"d7", -- 6290
         x"bc",  x"d6",  x"03",  x"03",  x"90",  x"d0",  x"e3",  x"d3", -- 6298
         x"bd",  x"d0",  x"1f",  x"d9",  x"fd",  x"d9",  x"59",  x"d5", -- 62A0
         x"6d",  x"d9",  x"70",  x"da",  x"76",  x"da",  x"d7",  x"da", -- 62A8
         x"ec",  x"da",  x"31",  x"d4",  x"44",  x"d4",  x"d5",  x"d6", -- 62B0
         x"2c",  x"d3",  x"56",  x"d1",  x"bf",  x"d3",  x"3b",  x"d3", -- 62B8
         x"4b",  x"d3",  x"5b",  x"d3",  x"89",  x"d3",  x"92",  x"d3", -- 62C0
         x"79",  x"11",  x"d8",  x"79",  x"6a",  x"d4",  x"7c",  x"98", -- 62C8
         x"d5",  x"7c",  x"f3",  x"d5",  x"7f",  x"28",  x"d9",  x"50", -- 62D0
         x"5e",  x"ce",  x"46",  x"5d",  x"ce",  x"4e",  x"46",  x"53", -- 62D8
         x"4e",  x"52",  x"47",  x"4f",  x"44",  x"46",  x"43",  x"4f", -- 62E0
         x"56",  x"4f",  x"4d",  x"55",  x"4c",  x"42",  x"53",  x"44", -- 62E8
         x"44",  x"2f",  x"30",  x"49",  x"44",  x"54",  x"4d",  x"4f", -- 62F0
         x"53",  x"4c",  x"53",  x"53",  x"54",  x"43",  x"4e",  x"55", -- 62F8
         x"46",  x"4d",  x"4f",  x"49",  x"4f",  x"20",  x"45",  x"52", -- 6300
         x"52",  x"4f",  x"52",  x"07",  x"00",  x"20",  x"49",  x"4e", -- 6308
         x"20",  x"00",  x"46",  x"49",  x"4c",  x"45",  x"20",  x"46", -- 6310
         x"4f",  x"55",  x"4e",  x"44",  x"0d",  x"4f",  x"4b",  x"0d", -- 6318
         x"00",  x"42",  x"52",  x"45",  x"41",  x"4b",  x"00",  x"e5", -- 6320
         x"2a",  x"db",  x"03",  x"06",  x"00",  x"09",  x"09",  x"3e", -- 6328
         x"e5",  x"3e",  x"d0",  x"95",  x"6f",  x"3e",  x"ff",  x"9c", -- 6330
         x"38",  x"04",  x"67",  x"39",  x"e1",  x"d8",  x"1e",  x"0c", -- 6338
         x"18",  x"14",  x"2a",  x"ca",  x"03",  x"22",  x"58",  x"03", -- 6340
         x"1e",  x"02",  x"01",  x"1e",  x"14",  x"01",  x"1e",  x"00", -- 6348
         x"01",  x"1e",  x"12",  x"01",  x"1e",  x"22",  x"cd",  x"69", -- 6350
         x"c6",  x"32",  x"43",  x"03",  x"cd",  x"55",  x"cb",  x"21", -- 6358
         x"dd",  x"c2",  x"57",  x"19",  x"44",  x"4d",  x"0b",  x"3e", -- 6360
         x"3f",  x"1e",  x"03",  x"cd",  x"d6",  x"d1",  x"21",  x"05", -- 6368
         x"c3",  x"cd",  x"c9",  x"d1",  x"2a",  x"58",  x"03",  x"11", -- 6370
         x"fe",  x"ff",  x"cd",  x"89",  x"c6",  x"ca",  x"0d",  x"c0", -- 6378
         x"7c",  x"a5",  x"3c",  x"c4",  x"21",  x"d8",  x"3e",  x"c1", -- 6380
         x"af",  x"32",  x"43",  x"03",  x"cd",  x"55",  x"cb",  x"21", -- 6388
         x"1d",  x"c3",  x"cd",  x"c9",  x"d1",  x"37",  x"dc",  x"fd", -- 6390
         x"dd",  x"cd",  x"df",  x"c6",  x"2b",  x"22",  x"58",  x"03", -- 6398
         x"21",  x"ea",  x"03",  x"3a",  x"4d",  x"03",  x"b7",  x"28", -- 63A0
         x"6b",  x"ed",  x"5b",  x"4e",  x"03",  x"f2",  x"f0",  x"c3", -- 63A8
         x"d5",  x"cd",  x"2a",  x"d8",  x"d1",  x"d5",  x"cd",  x"bb", -- 63B0
         x"c4",  x"3e",  x"2a",  x"38",  x"02",  x"3e",  x"20",  x"cd", -- 63B8
         x"ae",  x"c6",  x"cd",  x"ae",  x"c5",  x"d1",  x"30",  x"06", -- 63C0
         x"af",  x"32",  x"4d",  x"03",  x"18",  x"ba",  x"2a",  x"50", -- 63C8
         x"03",  x"19",  x"38",  x"f4",  x"d5",  x"11",  x"f9",  x"ff", -- 63D0
         x"cd",  x"89",  x"c6",  x"d1",  x"30",  x"ea",  x"22",  x"4e", -- 63D8
         x"03",  x"21",  x"62",  x"03",  x"f5",  x"18",  x"47",  x"c8", -- 63E0
         x"cd",  x"97",  x"c6",  x"cd",  x"86",  x"c9",  x"c0",  x"c1", -- 63E8
         x"cd",  x"bb",  x"c4",  x"30",  x"58",  x"d5",  x"7e",  x"23", -- 63F0
         x"b6",  x"23",  x"28",  x"02",  x"3e",  x"7f",  x"32",  x"4d", -- 63F8
         x"03",  x"7e",  x"23",  x"66",  x"6f",  x"22",  x"4e",  x"03", -- 6400
         x"cd",  x"98",  x"de",  x"d1",  x"c2",  x"96",  x"c3",  x"38", -- 6408
         x"b7",  x"3f",  x"18",  x"cd",  x"3e",  x"3e",  x"cd",  x"ae", -- 6410
         x"c6",  x"cd",  x"ae",  x"c5",  x"da",  x"96",  x"c3",  x"21", -- 6418
         x"61",  x"03",  x"cd",  x"bd",  x"c8",  x"3c",  x"3d",  x"ca", -- 6420
         x"96",  x"c3",  x"f5",  x"cd",  x"86",  x"c9",  x"d5",  x"cd", -- 6428
         x"da",  x"c4",  x"47",  x"d1",  x"f1",  x"d2",  x"8a",  x"c8", -- 6430
         x"d5",  x"c5",  x"af",  x"32",  x"cd",  x"03",  x"cd",  x"bd", -- 6438
         x"c8",  x"b7",  x"f5",  x"cd",  x"bb",  x"c4",  x"38",  x"08", -- 6440
         x"f1",  x"f5",  x"b7",  x"20",  x"03",  x"c3",  x"20",  x"ca", -- 6448
         x"c5",  x"30",  x"11",  x"eb",  x"2a",  x"d7",  x"03",  x"1a", -- 6450
         x"02",  x"03",  x"13",  x"cd",  x"89",  x"c6",  x"20",  x"f7", -- 6458
         x"ed",  x"43",  x"d7",  x"03",  x"d1",  x"f1",  x"28",  x"22", -- 6460
         x"2a",  x"d7",  x"03",  x"e3",  x"c1",  x"09",  x"e5",  x"cd", -- 6468
         x"ab",  x"c4",  x"e1",  x"22",  x"d7",  x"03",  x"eb",  x"36", -- 6470
         x"ff",  x"d1",  x"23",  x"23",  x"73",  x"23",  x"72",  x"23", -- 6478
         x"11",  x"62",  x"03",  x"1a",  x"77",  x"23",  x"13",  x"b7", -- 6480
         x"20",  x"f9",  x"cd",  x"4f",  x"c6",  x"23",  x"eb",  x"21", -- 6488
         x"96",  x"c3",  x"e5",  x"62",  x"6b",  x"7e",  x"23",  x"b6", -- 6490
         x"c8",  x"23",  x"7e",  x"23",  x"a6",  x"3c",  x"c8",  x"23", -- 6498
         x"af",  x"be",  x"23",  x"20",  x"fc",  x"eb",  x"73",  x"23", -- 64A0
         x"72",  x"18",  x"e8",  x"cd",  x"30",  x"c3",  x"c5",  x"e3", -- 64A8
         x"c1",  x"cd",  x"89",  x"c6",  x"7e",  x"02",  x"c8",  x"0b", -- 64B0
         x"2b",  x"18",  x"f6",  x"2a",  x"5f",  x"03",  x"44",  x"4d", -- 64B8
         x"7e",  x"23",  x"b6",  x"2b",  x"c8",  x"23",  x"23",  x"7e", -- 64C0
         x"23",  x"66",  x"6f",  x"cd",  x"89",  x"c6",  x"60",  x"69", -- 64C8
         x"7e",  x"23",  x"66",  x"6f",  x"3f",  x"c8",  x"3f",  x"d0", -- 64D0
         x"18",  x"e4",  x"af",  x"32",  x"af",  x"03",  x"0e",  x"05", -- 64D8
         x"11",  x"62",  x"03",  x"af",  x"32",  x"fb",  x"03",  x"7e", -- 64E0
         x"fe",  x"20",  x"ca",  x"71",  x"c5",  x"47",  x"fe",  x"22", -- 64E8
         x"ca",  x"91",  x"c5",  x"b7",  x"ca",  x"97",  x"c5",  x"3a", -- 64F0
         x"af",  x"03",  x"b7",  x"7e",  x"20",  x"73",  x"fe",  x"3f", -- 64F8
         x"3e",  x"9e",  x"28",  x"6d",  x"7e",  x"fe",  x"30",  x"38", -- 6500
         x"04",  x"fe",  x"3c",  x"38",  x"64",  x"d5",  x"11",  x"20", -- 6508
         x"c1",  x"c5",  x"01",  x"6d",  x"c5",  x"c5",  x"06",  x"7f", -- 6510
         x"7e",  x"fe",  x"61",  x"38",  x"07",  x"fe",  x"7b",  x"30", -- 6518
         x"03",  x"e6",  x"5f",  x"77",  x"4e",  x"eb",  x"23",  x"b6", -- 6520
         x"f2",  x"26",  x"c5",  x"04",  x"7e",  x"e6",  x"7f",  x"20", -- 6528
         x"15",  x"3a",  x"fc",  x"03",  x"a7",  x"c8",  x"3a",  x"fb", -- 6530
         x"03",  x"a7",  x"c0",  x"3c",  x"32",  x"fb",  x"03",  x"2a", -- 6538
         x"0c",  x"e0",  x"7e",  x"e6",  x"7f",  x"c8",  x"b9",  x"20", -- 6540
         x"dd",  x"eb",  x"e5",  x"13",  x"1a",  x"b7",  x"fa",  x"69", -- 6548
         x"c5",  x"4f",  x"78",  x"fe",  x"88",  x"20",  x"04",  x"cd", -- 6550
         x"bd",  x"c8",  x"2b",  x"23",  x"7e",  x"fe",  x"61",  x"38", -- 6558
         x"02",  x"e6",  x"5f",  x"b9",  x"28",  x"e5",  x"e1",  x"18", -- 6560
         x"bb",  x"48",  x"f1",  x"eb",  x"c9",  x"eb",  x"79",  x"c1", -- 6568
         x"d1",  x"23",  x"12",  x"13",  x"0c",  x"d6",  x"3a",  x"28", -- 6570
         x"04",  x"fe",  x"49",  x"20",  x"03",  x"32",  x"af",  x"03", -- 6578
         x"d6",  x"54",  x"28",  x"05",  x"d6",  x"0e",  x"c2",  x"e3", -- 6580
         x"c4",  x"47",  x"7e",  x"b7",  x"28",  x"09",  x"b8",  x"28", -- 6588
         x"e0",  x"23",  x"12",  x"0c",  x"13",  x"18",  x"f3",  x"21", -- 6590
         x"61",  x"03",  x"12",  x"13",  x"12",  x"13",  x"12",  x"c9", -- 6598
         x"4c",  x"49",  x"53",  x"54",  x"00",  x"52",  x"55",  x"4e", -- 65A0
         x"00",  x"43",  x"4f",  x"4e",  x"54",  x"00",  x"e5",  x"21", -- 65A8
         x"62",  x"03",  x"e3",  x"cd",  x"e4",  x"dd",  x"e3",  x"fe", -- 65B0
         x"1c",  x"11",  x"9f",  x"c5",  x"28",  x"0e",  x"fe",  x"1d", -- 65B8
         x"11",  x"a4",  x"c5",  x"28",  x"07",  x"fe",  x"1e",  x"11", -- 65C0
         x"a8",  x"c5",  x"20",  x"14",  x"21",  x"61",  x"03",  x"23", -- 65C8
         x"13",  x"1a",  x"77",  x"a7",  x"20",  x"f9",  x"21",  x"62", -- 65D0
         x"03",  x"cd",  x"f1",  x"c5",  x"e1",  x"c3",  x"5e",  x"cb", -- 65D8
         x"cd",  x"0f",  x"df",  x"20",  x"02",  x"e1",  x"c9",  x"cd", -- 65E0
         x"27",  x"df",  x"38",  x"f9",  x"cd",  x"32",  x"df",  x"18", -- 65E8
         x"c1",  x"7e",  x"b7",  x"c8",  x"cd",  x"d5",  x"dd",  x"23", -- 65F0
         x"18",  x"f7",  x"11",  x"0a",  x"00",  x"d5",  x"28",  x"17", -- 65F8
         x"cd",  x"86",  x"c9",  x"eb",  x"e3",  x"28",  x"11",  x"eb", -- 6600
         x"cd",  x"d6",  x"c8",  x"ed",  x"5b",  x"50",  x"03",  x"28", -- 6608
         x"06",  x"cd",  x"86",  x"c9",  x"c2",  x"48",  x"c3",  x"eb", -- 6610
         x"7d",  x"b4",  x"ca",  x"67",  x"c9",  x"22",  x"50",  x"03", -- 6618
         x"cb",  x"ff",  x"32",  x"4d",  x"03",  x"e1",  x"22",  x"4e", -- 6620
         x"03",  x"c1",  x"c3",  x"96",  x"c3",  x"cd",  x"5f",  x"de", -- 6628
         x"3a",  x"09",  x"03",  x"e6",  x"03",  x"28",  x"f3",  x"3e", -- 6630
         x"d5",  x"cd",  x"b2",  x"dc",  x"f1",  x"af",  x"18",  x"ea", -- 6638
         x"c0",  x"2a",  x"5f",  x"03",  x"af",  x"32",  x"5e",  x"03", -- 6640
         x"77",  x"23",  x"77",  x"23",  x"22",  x"d7",  x"03",  x"2a", -- 6648
         x"5f",  x"03",  x"2b",  x"22",  x"cf",  x"03",  x"2a",  x"b0", -- 6650
         x"03",  x"22",  x"c4",  x"03",  x"af",  x"cd",  x"df",  x"c8", -- 6658
         x"2a",  x"d7",  x"03",  x"22",  x"d9",  x"03",  x"22",  x"db", -- 6660
         x"03",  x"c1",  x"2a",  x"56",  x"03",  x"f9",  x"21",  x"b4", -- 6668
         x"03",  x"22",  x"b2",  x"03",  x"cd",  x"1d",  x"de",  x"af", -- 6670
         x"6f",  x"67",  x"22",  x"d5",  x"03",  x"32",  x"cc",  x"03", -- 6678
         x"22",  x"df",  x"03",  x"e5",  x"c5",  x"2a",  x"cf",  x"03", -- 6680
         x"c9",  x"7c",  x"92",  x"c0",  x"7d",  x"93",  x"c9",  x"7e", -- 6688
         x"fe",  x"41",  x"d8",  x"fe",  x"5b",  x"3f",  x"c9",  x"3a", -- 6690
         x"5e",  x"03",  x"a7",  x"c8",  x"cd",  x"69",  x"c6",  x"c3", -- 6698
         x"6e",  x"c3",  x"cd",  x"89",  x"c6",  x"3e",  x"08",  x"18", -- 66A0
         x"02",  x"3e",  x"20",  x"c3",  x"d5",  x"dd",  x"f5",  x"c5", -- 66A8
         x"4f",  x"fe",  x"20",  x"38",  x"13",  x"3a",  x"41",  x"03", -- 66B0
         x"47",  x"3a",  x"ac",  x"03",  x"04",  x"28",  x"05",  x"05", -- 66B8
         x"b8",  x"cc",  x"61",  x"cb",  x"3c",  x"32",  x"ac",  x"03", -- 66C0
         x"79",  x"cd",  x"d5",  x"dd",  x"c1",  x"f1",  x"c9",  x"3e", -- 66C8
         x"3f",  x"cd",  x"ae",  x"c6",  x"3e",  x"09",  x"cd",  x"ae", -- 66D0
         x"c6",  x"cd",  x"df",  x"c6",  x"c3",  x"4a",  x"03",  x"21", -- 66D8
         x"00",  x"20",  x"22",  x"61",  x"03",  x"22",  x"63",  x"03", -- 66E0
         x"65",  x"c9",  x"cd",  x"6c",  x"c9",  x"ed",  x"53",  x"46", -- 66E8
         x"03",  x"c9",  x"cd",  x"97",  x"c6",  x"cd",  x"25",  x"de", -- 66F0
         x"cd",  x"c8",  x"dd",  x"28",  x"12",  x"3e",  x"d5",  x"cd", -- 66F8
         x"b2",  x"dc",  x"2a",  x"46",  x"03",  x"22",  x"4e",  x"03", -- 6700
         x"21",  x"ff",  x"ff",  x"22",  x"46",  x"03",  x"e1",  x"cd", -- 6708
         x"86",  x"c9",  x"c0",  x"c1",  x"cd",  x"bb",  x"c4",  x"c5", -- 6710
         x"cd",  x"91",  x"c7",  x"e1",  x"4e",  x"23",  x"46",  x"23", -- 6718
         x"78",  x"b1",  x"28",  x"59",  x"cd",  x"67",  x"c7",  x"cd", -- 6720
         x"f9",  x"c8",  x"c5",  x"5e",  x"23",  x"56",  x"23",  x"e5", -- 6728
         x"21",  x"ea",  x"03",  x"cd",  x"61",  x"cb",  x"cd",  x"2a", -- 6730
         x"d8",  x"3e",  x"20",  x"e1",  x"cd",  x"ae",  x"c6",  x"7e", -- 6738
         x"23",  x"fe",  x"22",  x"28",  x"14",  x"b7",  x"28",  x"d3", -- 6740
         x"f2",  x"3c",  x"c7",  x"cd",  x"9a",  x"c7",  x"cd",  x"ae", -- 6748
         x"c6",  x"1a",  x"13",  x"b7",  x"f2",  x"4e",  x"c7",  x"18", -- 6750
         x"e6",  x"cd",  x"ae",  x"c6",  x"7e",  x"23",  x"b7",  x"28", -- 6758
         x"ba",  x"fe",  x"22",  x"28",  x"d7",  x"18",  x"f2",  x"e5", -- 6760
         x"2a",  x"44",  x"03",  x"7d",  x"b4",  x"2b",  x"22",  x"44", -- 6768
         x"03",  x"e1",  x"c0",  x"cd",  x"91",  x"c7",  x"cd",  x"e4", -- 6770
         x"dd",  x"fe",  x"03",  x"20",  x"ea",  x"cd",  x"c8",  x"dd", -- 6778
         x"28",  x"0c",  x"cd",  x"61",  x"cb",  x"cd",  x"fd",  x"dd", -- 6780
         x"2a",  x"4e",  x"03",  x"22",  x"46",  x"03",  x"c3",  x"8c", -- 6788
         x"c0",  x"e5",  x"2a",  x"46",  x"03",  x"22",  x"44",  x"03", -- 6790
         x"e1",  x"c9",  x"d6",  x"7f",  x"fe",  x"56",  x"38",  x"08", -- 6798
         x"d6",  x"55",  x"ed",  x"5b",  x"0c",  x"e0",  x"18",  x"03", -- 67A0
         x"11",  x"21",  x"c1",  x"47",  x"1a",  x"13",  x"b7",  x"f2", -- 67A8
         x"ac",  x"c7",  x"10",  x"f8",  x"e6",  x"7f",  x"c9",  x"3e", -- 67B0
         x"af",  x"32",  x"0a",  x"03",  x"c9",  x"21",  x"04",  x"00", -- 67B8
         x"39",  x"7e",  x"23",  x"fe",  x"81",  x"c0",  x"4e",  x"23", -- 67C0
         x"46",  x"23",  x"e5",  x"69",  x"60",  x"7a",  x"b3",  x"eb", -- 67C8
         x"28",  x"04",  x"eb",  x"cd",  x"89",  x"c6",  x"01",  x"0d", -- 67D0
         x"00",  x"e1",  x"c8",  x"09",  x"18",  x"e3",  x"3e",  x"64", -- 67D8
         x"32",  x"cc",  x"03",  x"cd",  x"5d",  x"ca",  x"c1",  x"e5", -- 67E0
         x"cd",  x"48",  x"ca",  x"22",  x"c8",  x"03",  x"21",  x"02", -- 67E8
         x"00",  x"39",  x"cd",  x"c1",  x"c7",  x"d1",  x"20",  x"14", -- 67F0
         x"09",  x"d5",  x"2b",  x"56",  x"2b",  x"5e",  x"23",  x"23", -- 67F8
         x"e5",  x"2a",  x"c8",  x"03",  x"cd",  x"89",  x"c6",  x"e1", -- 6800
         x"20",  x"e8",  x"d1",  x"f9",  x"eb",  x"0e",  x"08",  x"cd", -- 6808
         x"27",  x"c3",  x"e5",  x"2a",  x"c8",  x"03",  x"e3",  x"e5", -- 6810
         x"2a",  x"58",  x"03",  x"e3",  x"cd",  x"29",  x"cd",  x"cd", -- 6818
         x"cc",  x"c8",  x"a6",  x"cd",  x"26",  x"cd",  x"e5",  x"cd", -- 6820
         x"eb",  x"d6",  x"e1",  x"c5",  x"d5",  x"01",  x"00",  x"81", -- 6828
         x"51",  x"5a",  x"7e",  x"fe",  x"ab",  x"3e",  x"01",  x"20", -- 6830
         x"0e",  x"cd",  x"bd",  x"c8",  x"cd",  x"26",  x"cd",  x"e5", -- 6838
         x"cd",  x"eb",  x"d6",  x"cd",  x"97",  x"d6",  x"e1",  x"c5", -- 6840
         x"d5",  x"f5",  x"33",  x"e5",  x"2a",  x"cf",  x"03",  x"e3", -- 6848
         x"06",  x"81",  x"c5",  x"33",  x"cd",  x"16",  x"de",  x"cd", -- 6850
         x"f9",  x"c8",  x"22",  x"cf",  x"03",  x"7e",  x"fe",  x"3a", -- 6858
         x"28",  x"28",  x"b7",  x"c2",  x"48",  x"c3",  x"23",  x"7e", -- 6860
         x"23",  x"b6",  x"ca",  x"22",  x"c9",  x"23",  x"5e",  x"23", -- 6868
         x"56",  x"ed",  x"53",  x"58",  x"03",  x"3a",  x"0a",  x"03", -- 6870
         x"b7",  x"28",  x"0f",  x"e5",  x"3e",  x"3c",  x"cd",  x"ae", -- 6878
         x"c6",  x"cd",  x"2a",  x"d8",  x"3e",  x"3e",  x"cd",  x"ae", -- 6880
         x"c6",  x"e1",  x"cd",  x"bd",  x"c8",  x"11",  x"54",  x"c8", -- 6888
         x"d5",  x"c8",  x"d6",  x"80",  x"da",  x"5d",  x"ca",  x"fe", -- 6890
         x"25",  x"38",  x"14",  x"d6",  x"50",  x"38",  x"34",  x"fe", -- 6898
         x"05",  x"38",  x"0a",  x"47",  x"3a",  x"fc",  x"03",  x"a7", -- 68A0
         x"28",  x"29",  x"c3",  x"03",  x"e0",  x"c6",  x"25",  x"07", -- 68A8
         x"4f",  x"06",  x"00",  x"eb",  x"21",  x"40",  x"c2",  x"09", -- 68B0
         x"4e",  x"23",  x"46",  x"c5",  x"eb",  x"23",  x"7e",  x"fe", -- 68B8
         x"3a",  x"d0",  x"fe",  x"20",  x"28",  x"f7",  x"fe",  x"30", -- 68C0
         x"3f",  x"3c",  x"3d",  x"c9",  x"7e",  x"e3",  x"be",  x"23", -- 68C8
         x"e3",  x"28",  x"ea",  x"c3",  x"48",  x"c3",  x"3e",  x"2c", -- 68D0
         x"be",  x"18",  x"f6",  x"3e",  x"29",  x"18",  x"f9",  x"eb", -- 68D8
         x"2a",  x"5f",  x"03",  x"28",  x"0e",  x"eb",  x"cd",  x"86", -- 68E0
         x"c9",  x"e5",  x"cd",  x"bb",  x"c4",  x"60",  x"69",  x"d1", -- 68E8
         x"d2",  x"20",  x"ca",  x"2b",  x"22",  x"dd",  x"03",  x"eb", -- 68F0
         x"c9",  x"cd",  x"f3",  x"dd",  x"c0",  x"fe",  x"13",  x"28", -- 68F8
         x"08",  x"fe",  x"03",  x"c0",  x"cd",  x"e4",  x"dd",  x"18", -- 6900
         x"0f",  x"cd",  x"e4",  x"dd",  x"fe",  x"1e",  x"c8",  x"fe", -- 6908
         x"0a",  x"c8",  x"fe",  x"03",  x"28",  x"02",  x"18",  x"f1", -- 6910
         x"c0",  x"f6",  x"c0",  x"22",  x"cf",  x"03",  x"21",  x"f6", -- 6918
         x"ff",  x"c1",  x"2a",  x"58",  x"03",  x"f5",  x"7d",  x"a4", -- 6920
         x"3c",  x"28",  x"09",  x"22",  x"d3",  x"03",  x"2a",  x"cf", -- 6928
         x"03",  x"22",  x"d5",  x"03",  x"af",  x"32",  x"43",  x"03", -- 6930
         x"cd",  x"1d",  x"de",  x"cd",  x"55",  x"cb",  x"f1",  x"21", -- 6938
         x"21",  x"c3",  x"c2",  x"71",  x"c3",  x"c3",  x"88",  x"c3", -- 6940
         x"2a",  x"d5",  x"03",  x"7c",  x"b5",  x"1e",  x"20",  x"ca", -- 6948
         x"56",  x"c3",  x"eb",  x"2a",  x"d3",  x"03",  x"22",  x"58", -- 6950
         x"03",  x"eb",  x"c9",  x"cd",  x"bd",  x"c8",  x"cd",  x"26", -- 6958
         x"cd",  x"cd",  x"97",  x"d6",  x"f2",  x"6f",  x"c9",  x"1e", -- 6960
         x"08",  x"c3",  x"56",  x"c3",  x"cd",  x"26",  x"cd",  x"3a", -- 6968
         x"e8",  x"03",  x"fe",  x"90",  x"da",  x"45",  x"d7",  x"01", -- 6970
         x"80",  x"90",  x"11",  x"00",  x"00",  x"e5",  x"cd",  x"18", -- 6978
         x"d7",  x"e1",  x"51",  x"c8",  x"18",  x"e1",  x"2b",  x"11", -- 6980
         x"00",  x"00",  x"cd",  x"bd",  x"c8",  x"d0",  x"e5",  x"f5", -- 6988
         x"21",  x"98",  x"19",  x"cd",  x"89",  x"c6",  x"da",  x"48", -- 6990
         x"c3",  x"62",  x"6b",  x"19",  x"29",  x"19",  x"29",  x"f1", -- 6998
         x"d6",  x"30",  x"5f",  x"16",  x"00",  x"19",  x"eb",  x"e1", -- 69A0
         x"18",  x"e0",  x"28",  x"3c",  x"cd",  x"5e",  x"c9",  x"cd", -- 69A8
         x"be",  x"c8",  x"e5",  x"2a",  x"b0",  x"03",  x"28",  x"10", -- 69B0
         x"e1",  x"cd",  x"d6",  x"c8",  x"d5",  x"cd",  x"6c",  x"c9", -- 69B8
         x"cd",  x"be",  x"c8",  x"c2",  x"48",  x"c3",  x"e3",  x"eb", -- 69C0
         x"7d",  x"93",  x"5f",  x"7c",  x"9a",  x"57",  x"da",  x"3e", -- 69C8
         x"c3",  x"e5",  x"2a",  x"d7",  x"03",  x"01",  x"28",  x"00", -- 69D0
         x"09",  x"cd",  x"89",  x"c6",  x"d2",  x"3e",  x"c3",  x"eb", -- 69D8
         x"22",  x"56",  x"03",  x"e1",  x"22",  x"b0",  x"03",  x"e1", -- 69E0
         x"c3",  x"53",  x"c6",  x"ca",  x"4f",  x"c6",  x"cd",  x"53", -- 69E8
         x"c6",  x"01",  x"54",  x"c8",  x"18",  x"10",  x"0e",  x"03", -- 69F0
         x"cd",  x"27",  x"c3",  x"c1",  x"e5",  x"e5",  x"2a",  x"58", -- 69F8
         x"03",  x"e3",  x"3e",  x"8c",  x"f5",  x"33",  x"c5",  x"cd", -- 6A00
         x"86",  x"c9",  x"cd",  x"4a",  x"ca",  x"e5",  x"2a",  x"58", -- 6A08
         x"03",  x"cd",  x"89",  x"c6",  x"e1",  x"23",  x"dc",  x"be", -- 6A10
         x"c4",  x"d4",  x"bb",  x"c4",  x"60",  x"69",  x"2b",  x"d8", -- 6A18
         x"1e",  x"0e",  x"c3",  x"56",  x"c3",  x"c0",  x"16",  x"ff", -- 6A20
         x"cd",  x"bd",  x"c7",  x"f9",  x"fe",  x"8c",  x"1e",  x"04", -- 6A28
         x"20",  x"f0",  x"e1",  x"22",  x"58",  x"03",  x"23",  x"7c", -- 6A30
         x"b5",  x"20",  x"07",  x"3a",  x"cd",  x"03",  x"b7",  x"c2", -- 6A38
         x"87",  x"c3",  x"21",  x"54",  x"c8",  x"e3",  x"3e",  x"e1", -- 6A40
         x"01",  x"3a",  x"0e",  x"00",  x"06",  x"00",  x"79",  x"48", -- 6A48
         x"47",  x"7e",  x"b7",  x"c8",  x"b8",  x"c8",  x"23",  x"fe", -- 6A50
         x"22",  x"28",  x"f3",  x"18",  x"f4",  x"cd",  x"06",  x"cf", -- 6A58
         x"cd",  x"cc",  x"c8",  x"b4",  x"d5",  x"3a",  x"ae",  x"03", -- 6A60
         x"f5",  x"cd",  x"3a",  x"cd",  x"f1",  x"e3",  x"22",  x"cf", -- 6A68
         x"03",  x"1f",  x"cd",  x"2b",  x"cd",  x"28",  x"35",  x"e5", -- 6A70
         x"2a",  x"e5",  x"03",  x"e5",  x"23",  x"23",  x"5e",  x"23", -- 6A78
         x"56",  x"2a",  x"5f",  x"03",  x"cd",  x"89",  x"c6",  x"30", -- 6A80
         x"12",  x"2a",  x"56",  x"03",  x"cd",  x"89",  x"c6",  x"d1", -- 6A88
         x"30",  x"11",  x"21",  x"c0",  x"03",  x"cd",  x"89",  x"c6", -- 6A90
         x"30",  x"09",  x"3e",  x"d1",  x"cd",  x"1b",  x"d3",  x"eb", -- 6A98
         x"cd",  x"66",  x"d1",  x"cd",  x"1b",  x"d3",  x"e1",  x"cd", -- 6AA0
         x"fa",  x"d6",  x"e1",  x"c9",  x"e5",  x"cd",  x"f7",  x"d6", -- 6AA8
         x"d1",  x"e1",  x"c9",  x"cd",  x"21",  x"d4",  x"7e",  x"47", -- 6AB0
         x"fe",  x"8c",  x"28",  x"05",  x"cd",  x"cc",  x"c8",  x"88", -- 6AB8
         x"2b",  x"4b",  x"0d",  x"78",  x"ca",  x"92",  x"c8",  x"cd", -- 6AC0
         x"87",  x"c9",  x"fe",  x"2c",  x"c0",  x"18",  x"f3",  x"cd", -- 6AC8
         x"3a",  x"cd",  x"7e",  x"fe",  x"88",  x"28",  x"05",  x"cd", -- 6AD0
         x"cc",  x"c8",  x"a9",  x"2b",  x"cd",  x"29",  x"cd",  x"cd", -- 6AD8
         x"97",  x"d6",  x"20",  x"08",  x"23",  x"7e",  x"b7",  x"c8", -- 6AE0
         x"fe",  x"d4",  x"20",  x"f8",  x"cd",  x"bd",  x"c8",  x"da", -- 6AE8
         x"07",  x"ca",  x"c3",  x"91",  x"c8",  x"cd",  x"be",  x"c8", -- 6AF0
         x"18",  x"07",  x"af",  x"32",  x"fd",  x"03",  x"cd",  x"25", -- 6AF8
         x"de",  x"28",  x"5e",  x"c8",  x"fe",  x"d5",  x"38",  x"09", -- 6B00
         x"3a",  x"fc",  x"03",  x"a7",  x"28",  x"03",  x"cd",  x"06", -- 6B08
         x"e0",  x"fe",  x"a5",  x"ca",  x"92",  x"cb",  x"fe",  x"a8", -- 6B10
         x"28",  x"78",  x"e5",  x"fe",  x"2c",  x"28",  x"5d",  x"fe", -- 6B18
         x"3b",  x"ca",  x"b2",  x"cb",  x"c1",  x"cd",  x"3a",  x"cd", -- 6B20
         x"e5",  x"3a",  x"ae",  x"03",  x"b7",  x"20",  x"20",  x"cd", -- 6B28
         x"34",  x"d8",  x"cd",  x"8a",  x"d1",  x"36",  x"20",  x"2a", -- 6B30
         x"e5",  x"03",  x"34",  x"2a",  x"e5",  x"03",  x"3a",  x"41", -- 6B38
         x"03",  x"47",  x"04",  x"28",  x"0a",  x"04",  x"3a",  x"ac", -- 6B40
         x"03",  x"86",  x"3d",  x"b8",  x"d4",  x"61",  x"cb",  x"cd", -- 6B48
         x"cc",  x"d1",  x"e1",  x"18",  x"a0",  x"3a",  x"ac",  x"03", -- 6B50
         x"b7",  x"c8",  x"18",  x"05",  x"36",  x"00",  x"21",  x"61", -- 6B58
         x"03",  x"3e",  x"0d",  x"cd",  x"ae",  x"c6",  x"3e",  x"0a", -- 6B60
         x"cd",  x"ae",  x"c6",  x"af",  x"32",  x"ac",  x"03",  x"3a", -- 6B68
         x"40",  x"03",  x"3d",  x"c8",  x"f5",  x"af",  x"cd",  x"ae", -- 6B70
         x"c6",  x"f1",  x"18",  x"f6",  x"3a",  x"42",  x"03",  x"47", -- 6B78
         x"3a",  x"ac",  x"03",  x"b8",  x"d4",  x"61",  x"cb",  x"30", -- 6B80
         x"29",  x"d6",  x"0d",  x"38",  x"02",  x"20",  x"fa",  x"2f", -- 6B88
         x"18",  x"15",  x"f5",  x"cd",  x"1e",  x"d4",  x"cd",  x"db", -- 6B90
         x"c8",  x"2b",  x"f1",  x"d6",  x"a8",  x"e5",  x"28",  x"03", -- 6B98
         x"3a",  x"ac",  x"03",  x"2f",  x"83",  x"30",  x"0b",  x"3c", -- 6BA0
         x"28",  x"08",  x"47",  x"3e",  x"20",  x"cd",  x"ae",  x"c6", -- 6BA8
         x"10",  x"fb",  x"e1",  x"cd",  x"bd",  x"c8",  x"c3",  x"03", -- 6BB0
         x"cb",  x"cd",  x"21",  x"d4",  x"32",  x"41",  x"03",  x"c9", -- 6BB8
         x"cd",  x"21",  x"d4",  x"c0",  x"3c",  x"32",  x"40",  x"03", -- 6BC0
         x"c9",  x"3f",  x"52",  x"45",  x"44",  x"4f",  x"20",  x"46", -- 6BC8
         x"52",  x"4f",  x"4d",  x"20",  x"53",  x"54",  x"41",  x"52", -- 6BD0
         x"54",  x"0d",  x"00",  x"3a",  x"ce",  x"03",  x"b7",  x"c2", -- 6BD8
         x"42",  x"c3",  x"c1",  x"21",  x"c9",  x"cb",  x"cd",  x"c9", -- 6BE0
         x"d1",  x"c3",  x"85",  x"c6",  x"cd",  x"37",  x"d1",  x"cd", -- 6BE8
         x"5f",  x"de",  x"af",  x"32",  x"43",  x"03",  x"7e",  x"fe", -- 6BF0
         x"22",  x"20",  x"10",  x"cd",  x"8b",  x"d1",  x"cd",  x"cc", -- 6BF8
         x"c8",  x"3b",  x"e5",  x"cd",  x"cc",  x"d1",  x"cd",  x"d4", -- 6C00
         x"c6",  x"18",  x"04",  x"e5",  x"cd",  x"cf",  x"c6",  x"c1", -- 6C08
         x"38",  x"36",  x"21",  x"62",  x"03",  x"7e",  x"b7",  x"2b", -- 6C10
         x"c5",  x"28",  x"37",  x"36",  x"2c",  x"18",  x"05",  x"e5", -- 6C18
         x"2a",  x"dd",  x"03",  x"f6",  x"af",  x"32",  x"ce",  x"03", -- 6C20
         x"e3",  x"18",  x"03",  x"cd",  x"d6",  x"c8",  x"cd",  x"06", -- 6C28
         x"cf",  x"e3",  x"d5",  x"7e",  x"fe",  x"2c",  x"28",  x"1e", -- 6C30
         x"3a",  x"ce",  x"03",  x"b7",  x"20",  x"7d",  x"3e",  x"3f", -- 6C38
         x"cd",  x"ae",  x"c6",  x"cd",  x"cf",  x"c6",  x"d1",  x"c1", -- 6C40
         x"da",  x"1f",  x"c9",  x"21",  x"62",  x"03",  x"7e",  x"b7", -- 6C48
         x"2b",  x"c5",  x"ca",  x"47",  x"ca",  x"d5",  x"3a",  x"ae", -- 6C50
         x"03",  x"b7",  x"28",  x"21",  x"cd",  x"bd",  x"c8",  x"57", -- 6C58
         x"47",  x"fe",  x"22",  x"28",  x"0c",  x"3a",  x"ce",  x"03", -- 6C60
         x"b7",  x"57",  x"28",  x"02",  x"16",  x"3a",  x"06",  x"2c", -- 6C68
         x"2b",  x"cd",  x"8e",  x"d1",  x"eb",  x"21",  x"88",  x"cc", -- 6C70
         x"e3",  x"d5",  x"c3",  x"77",  x"ca",  x"cd",  x"bd",  x"c8", -- 6C78
         x"cd",  x"a1",  x"d7",  x"e3",  x"cd",  x"f7",  x"d6",  x"e1", -- 6C80
         x"cd",  x"be",  x"c8",  x"28",  x"05",  x"fe",  x"2c",  x"c2", -- 6C88
         x"db",  x"cb",  x"e3",  x"cd",  x"be",  x"c8",  x"20",  x"93", -- 6C90
         x"d1",  x"3a",  x"ce",  x"03",  x"b7",  x"eb",  x"c2",  x"f4", -- 6C98
         x"c8",  x"d5",  x"b6",  x"21",  x"ab",  x"cc",  x"c4",  x"c9", -- 6CA0
         x"d1",  x"e1",  x"c9",  x"3f",  x"45",  x"58",  x"54",  x"52", -- 6CA8
         x"41",  x"20",  x"49",  x"47",  x"4e",  x"4f",  x"52",  x"45", -- 6CB0
         x"44",  x"0d",  x"00",  x"cd",  x"48",  x"ca",  x"b7",  x"20", -- 6CB8
         x"11",  x"23",  x"7e",  x"23",  x"b6",  x"1e",  x"06",  x"ca", -- 6CC0
         x"56",  x"c3",  x"23",  x"5e",  x"23",  x"56",  x"ed",  x"53", -- 6CC8
         x"ca",  x"03",  x"cd",  x"bd",  x"c8",  x"fe",  x"83",  x"20", -- 6CD0
         x"e2",  x"c3",  x"56",  x"cc",  x"11",  x"00",  x"00",  x"c4", -- 6CD8
         x"06",  x"cf",  x"22",  x"cf",  x"03",  x"cd",  x"bd",  x"c7", -- 6CE0
         x"c2",  x"4e",  x"c3",  x"f9",  x"d5",  x"7e",  x"23",  x"f5", -- 6CE8
         x"d5",  x"cd",  x"dd",  x"d6",  x"e3",  x"e5",  x"cd",  x"61", -- 6CF0
         x"d4",  x"e1",  x"cd",  x"f7",  x"d6",  x"e1",  x"cd",  x"ee", -- 6CF8
         x"d6",  x"e5",  x"cd",  x"18",  x"d7",  x"e1",  x"c1",  x"90", -- 6D00
         x"cd",  x"ee",  x"d6",  x"28",  x"09",  x"ed",  x"53",  x"58", -- 6D08
         x"03",  x"69",  x"60",  x"c3",  x"50",  x"c8",  x"f9",  x"2a", -- 6D10
         x"cf",  x"03",  x"7e",  x"fe",  x"2c",  x"c2",  x"54",  x"c8", -- 6D18
         x"cd",  x"bd",  x"c8",  x"cd",  x"df",  x"cc",  x"cd",  x"3a", -- 6D20
         x"cd",  x"f6",  x"37",  x"3a",  x"ae",  x"03",  x"8f",  x"b7", -- 6D28
         x"e8",  x"1e",  x"18",  x"c3",  x"56",  x"c3",  x"cd",  x"cc", -- 6D30
         x"c8",  x"28",  x"2b",  x"16",  x"00",  x"d5",  x"0e",  x"01", -- 6D38
         x"cd",  x"27",  x"c3",  x"cd",  x"ad",  x"cd",  x"22",  x"d1", -- 6D40
         x"03",  x"2a",  x"d1",  x"03",  x"c1",  x"78",  x"fe",  x"78", -- 6D48
         x"d4",  x"29",  x"cd",  x"7e",  x"16",  x"00",  x"d6",  x"b3", -- 6D50
         x"38",  x"15",  x"fe",  x"03",  x"30",  x"11",  x"fe",  x"01", -- 6D58
         x"17",  x"aa",  x"ba",  x"57",  x"da",  x"48",  x"c3",  x"22", -- 6D60
         x"c6",  x"03",  x"cd",  x"bd",  x"c8",  x"18",  x"e7",  x"7a", -- 6D68
         x"b7",  x"c2",  x"84",  x"ce",  x"7e",  x"22",  x"c6",  x"03", -- 6D70
         x"d6",  x"ac",  x"d8",  x"fe",  x"07",  x"d0",  x"5f",  x"3a", -- 6D78
         x"ae",  x"03",  x"3d",  x"b3",  x"7b",  x"ca",  x"b3",  x"d2", -- 6D80
         x"07",  x"83",  x"5f",  x"21",  x"c8",  x"c2",  x"19",  x"78", -- 6D88
         x"56",  x"ba",  x"d0",  x"23",  x"cd",  x"29",  x"cd",  x"c5", -- 6D90
         x"01",  x"49",  x"cd",  x"c5",  x"43",  x"4a",  x"cd",  x"c8", -- 6D98
         x"d6",  x"58",  x"51",  x"4e",  x"23",  x"46",  x"23",  x"c5", -- 6DA0
         x"2a",  x"c6",  x"03",  x"18",  x"90",  x"af",  x"32",  x"ae", -- 6DA8
         x"03",  x"cd",  x"bd",  x"c8",  x"1e",  x"24",  x"ca",  x"56", -- 6DB0
         x"c3",  x"da",  x"a1",  x"d7",  x"cd",  x"8f",  x"c6",  x"30", -- 6DB8
         x"37",  x"fe",  x"ac",  x"28",  x"e8",  x"fe",  x"2e",  x"ca", -- 6DC0
         x"a1",  x"d7",  x"fe",  x"ad",  x"28",  x"19",  x"fe",  x"22", -- 6DC8
         x"ca",  x"8b",  x"d1",  x"fe",  x"aa",  x"ca",  x"e3",  x"ce", -- 6DD0
         x"fe",  x"a7",  x"ca",  x"f0",  x"d0",  x"d6",  x"b6",  x"30", -- 6DD8
         x"28",  x"cd",  x"36",  x"cd",  x"c3",  x"db",  x"c8",  x"16", -- 6DE0
         x"7d",  x"cd",  x"3d",  x"cd",  x"2a",  x"d1",  x"03",  x"e5", -- 6DE8
         x"cd",  x"c0",  x"d6",  x"cd",  x"29",  x"cd",  x"e1",  x"c9", -- 6DF0
         x"cd",  x"06",  x"cf",  x"e5",  x"eb",  x"22",  x"e5",  x"03", -- 6DF8
         x"3a",  x"ae",  x"03",  x"b7",  x"cc",  x"dd",  x"d6",  x"e1", -- 6E00
         x"c9",  x"06",  x"00",  x"07",  x"4f",  x"c5",  x"cd",  x"bd", -- 6E08
         x"c8",  x"79",  x"fe",  x"33",  x"38",  x"07",  x"3a",  x"fc", -- 6E10
         x"03",  x"a7",  x"c2",  x"09",  x"e0",  x"fe",  x"22",  x"28", -- 6E18
         x"1e",  x"fe",  x"2d",  x"38",  x"17",  x"cd",  x"36",  x"cd", -- 6E20
         x"cd",  x"d6",  x"c8",  x"cd",  x"2a",  x"cd",  x"eb",  x"2a", -- 6E28
         x"e5",  x"03",  x"e3",  x"e5",  x"eb",  x"cd",  x"21",  x"d4", -- 6E30
         x"eb",  x"e3",  x"18",  x"08",  x"cd",  x"e1",  x"cd",  x"e3", -- 6E38
         x"11",  x"f3",  x"cd",  x"d5",  x"01",  x"94",  x"c2",  x"09", -- 6E40
         x"4e",  x"23",  x"66",  x"69",  x"e9",  x"15",  x"fe",  x"ad", -- 6E48
         x"c8",  x"fe",  x"2d",  x"c8",  x"14",  x"fe",  x"2b",  x"c8", -- 6E50
         x"fe",  x"ac",  x"c8",  x"2b",  x"c9",  x"f6",  x"af",  x"f5", -- 6E58
         x"cd",  x"29",  x"cd",  x"cd",  x"6f",  x"c9",  x"f1",  x"eb", -- 6E60
         x"c1",  x"e3",  x"eb",  x"cd",  x"e0",  x"d6",  x"f5",  x"cd", -- 6E68
         x"6f",  x"c9",  x"f1",  x"c1",  x"79",  x"21",  x"b0",  x"d0", -- 6E70
         x"20",  x"05",  x"a3",  x"4f",  x"78",  x"a2",  x"e9",  x"b3", -- 6E78
         x"4f",  x"78",  x"b2",  x"e9",  x"21",  x"96",  x"ce",  x"3a", -- 6E80
         x"ae",  x"03",  x"1f",  x"7a",  x"17",  x"5f",  x"16",  x"64", -- 6E88
         x"78",  x"ba",  x"d0",  x"c3",  x"97",  x"cd",  x"98",  x"ce", -- 6E90
         x"79",  x"b7",  x"1f",  x"c1",  x"d1",  x"f5",  x"cd",  x"2b", -- 6E98
         x"cd",  x"21",  x"d9",  x"ce",  x"e5",  x"ca",  x"18",  x"d7", -- 6EA0
         x"af",  x"32",  x"ae",  x"03",  x"d5",  x"cd",  x"fe",  x"d2", -- 6EA8
         x"7e",  x"23",  x"23",  x"4e",  x"23",  x"46",  x"d1",  x"c5", -- 6EB0
         x"f5",  x"cd",  x"02",  x"d3",  x"cd",  x"ee",  x"d6",  x"f1", -- 6EB8
         x"57",  x"e1",  x"7b",  x"b2",  x"c8",  x"7a",  x"d6",  x"01", -- 6EC0
         x"d8",  x"af",  x"bb",  x"3c",  x"d0",  x"15",  x"1d",  x"0a", -- 6EC8
         x"be",  x"23",  x"03",  x"28",  x"ed",  x"3f",  x"c3",  x"a2", -- 6ED0
         x"d6",  x"3c",  x"8f",  x"c1",  x"a0",  x"c6",  x"ff",  x"9f", -- 6ED8
         x"c3",  x"a9",  x"d6",  x"16",  x"5a",  x"cd",  x"3d",  x"cd", -- 6EE0
         x"cd",  x"29",  x"cd",  x"cd",  x"6f",  x"c9",  x"7b",  x"2f", -- 6EE8
         x"4f",  x"7a",  x"2f",  x"cd",  x"b0",  x"d0",  x"c1",  x"c3", -- 6EF0
         x"49",  x"cd",  x"cd",  x"be",  x"c8",  x"c8",  x"cd",  x"d6", -- 6EF8
         x"c8",  x"01",  x"fa",  x"ce",  x"c5",  x"f6",  x"af",  x"32", -- 6F00
         x"ad",  x"03",  x"46",  x"cd",  x"8f",  x"c6",  x"da",  x"48", -- 6F08
         x"c3",  x"af",  x"4f",  x"32",  x"ae",  x"03",  x"cd",  x"bd", -- 6F10
         x"c8",  x"38",  x"05",  x"cd",  x"8f",  x"c6",  x"38",  x"0b", -- 6F18
         x"4f",  x"cd",  x"bd",  x"c8",  x"38",  x"fb",  x"cd",  x"8f", -- 6F20
         x"c6",  x"30",  x"f6",  x"d6",  x"24",  x"20",  x"0a",  x"3c", -- 6F28
         x"32",  x"ae",  x"03",  x"0f",  x"81",  x"4f",  x"cd",  x"bd", -- 6F30
         x"c8",  x"3a",  x"cc",  x"03",  x"3d",  x"ca",  x"dd",  x"cf", -- 6F38
         x"f2",  x"48",  x"cf",  x"7e",  x"d6",  x"28",  x"28",  x"6f", -- 6F40
         x"af",  x"32",  x"cc",  x"03",  x"e5",  x"50",  x"59",  x"2a", -- 6F48
         x"df",  x"03",  x"cd",  x"89",  x"c6",  x"11",  x"e1",  x"03", -- 6F50
         x"ca",  x"e0",  x"d5",  x"2a",  x"d9",  x"03",  x"eb",  x"2a", -- 6F58
         x"d7",  x"03",  x"cd",  x"89",  x"c6",  x"28",  x"10",  x"79", -- 6F60
         x"96",  x"23",  x"20",  x"02",  x"78",  x"96",  x"23",  x"28", -- 6F68
         x"38",  x"23",  x"23",  x"23",  x"23",  x"18",  x"eb",  x"e1", -- 6F70
         x"e3",  x"d5",  x"11",  x"fb",  x"cd",  x"cd",  x"89",  x"c6", -- 6F78
         x"d1",  x"28",  x"29",  x"e3",  x"e5",  x"c5",  x"01",  x"06", -- 6F80
         x"00",  x"2a",  x"db",  x"03",  x"e5",  x"09",  x"c1",  x"e5", -- 6F88
         x"cd",  x"ab",  x"c4",  x"e1",  x"22",  x"db",  x"03",  x"60", -- 6F90
         x"69",  x"22",  x"d9",  x"03",  x"2b",  x"36",  x"00",  x"cd", -- 6F98
         x"89",  x"c6",  x"20",  x"f8",  x"d1",  x"73",  x"23",  x"72", -- 6FA0
         x"23",  x"eb",  x"e1",  x"c9",  x"32",  x"e8",  x"03",  x"21", -- 6FA8
         x"20",  x"c3",  x"22",  x"e5",  x"03",  x"e1",  x"c9",  x"e5", -- 6FB0
         x"2a",  x"ad",  x"03",  x"e3",  x"57",  x"d5",  x"c5",  x"cd", -- 6FB8
         x"5b",  x"c9",  x"c1",  x"f1",  x"eb",  x"e3",  x"e5",  x"eb", -- 6FC0
         x"3c",  x"57",  x"7e",  x"fe",  x"2c",  x"28",  x"ee",  x"cd", -- 6FC8
         x"db",  x"c8",  x"22",  x"d1",  x"03",  x"e1",  x"22",  x"ad", -- 6FD0
         x"03",  x"1e",  x"00",  x"d5",  x"11",  x"e5",  x"f5",  x"2a", -- 6FD8
         x"d9",  x"03",  x"3e",  x"19",  x"ed",  x"5b",  x"db",  x"03", -- 6FE0
         x"cd",  x"89",  x"c6",  x"28",  x"23",  x"7e",  x"b9",  x"23", -- 6FE8
         x"20",  x"02",  x"7e",  x"b8",  x"23",  x"5e",  x"23",  x"56", -- 6FF0
         x"23",  x"20",  x"e8",  x"3a",  x"ad",  x"03",  x"b7",  x"c2", -- 6FF8
         x"51",  x"c3",  x"f1",  x"44",  x"4d",  x"ca",  x"aa",  x"cf", -- 7000
         x"96",  x"28",  x"5f",  x"1e",  x"10",  x"c3",  x"56",  x"c3", -- 7008
         x"11",  x"04",  x"00",  x"f1",  x"ca",  x"67",  x"c9",  x"71", -- 7010
         x"23",  x"70",  x"23",  x"4f",  x"cd",  x"27",  x"c3",  x"23", -- 7018
         x"23",  x"22",  x"c6",  x"03",  x"71",  x"23",  x"3a",  x"ad", -- 7020
         x"03",  x"17",  x"79",  x"01",  x"0b",  x"00",  x"30",  x"02", -- 7028
         x"c1",  x"03",  x"71",  x"23",  x"70",  x"23",  x"f5",  x"e5", -- 7030
         x"cd",  x"89",  x"d7",  x"eb",  x"e1",  x"f1",  x"3d",  x"20", -- 7038
         x"ea",  x"f5",  x"42",  x"4b",  x"eb",  x"19",  x"da",  x"3e", -- 7040
         x"c3",  x"cd",  x"30",  x"c3",  x"22",  x"db",  x"03",  x"2b", -- 7048
         x"36",  x"00",  x"cd",  x"89",  x"c6",  x"20",  x"f8",  x"03", -- 7050
         x"57",  x"2a",  x"c6",  x"03",  x"5e",  x"eb",  x"29",  x"09", -- 7058
         x"eb",  x"2b",  x"2b",  x"73",  x"23",  x"72",  x"23",  x"f1", -- 7060
         x"38",  x"22",  x"47",  x"4f",  x"7e",  x"23",  x"16",  x"e1", -- 7068
         x"5e",  x"23",  x"56",  x"23",  x"e3",  x"f5",  x"cd",  x"89", -- 7070
         x"c6",  x"30",  x"90",  x"e5",  x"cd",  x"89",  x"d7",  x"d1", -- 7078
         x"19",  x"f1",  x"3d",  x"44",  x"4d",  x"20",  x"e8",  x"29", -- 7080
         x"29",  x"c1",  x"09",  x"eb",  x"2a",  x"d1",  x"03",  x"c9", -- 7088
         x"ed",  x"5b",  x"db",  x"03",  x"21",  x"00",  x"00",  x"39", -- 7090
         x"3a",  x"ae",  x"03",  x"b7",  x"28",  x"0d",  x"cd",  x"fe", -- 7098
         x"d2",  x"cd",  x"09",  x"d2",  x"ed",  x"5b",  x"56",  x"03", -- 70A0
         x"2a",  x"c4",  x"03",  x"7d",  x"93",  x"4f",  x"7c",  x"9a", -- 70A8
         x"41",  x"50",  x"1e",  x"00",  x"21",  x"ae",  x"03",  x"73", -- 70B0
         x"06",  x"90",  x"c3",  x"ae",  x"d6",  x"3a",  x"ac",  x"03", -- 70B8
         x"47",  x"af",  x"18",  x"ed",  x"cd",  x"45",  x"d1",  x"cd", -- 70C0
         x"37",  x"d1",  x"01",  x"48",  x"ca",  x"c5",  x"d5",  x"cd", -- 70C8
         x"cc",  x"c8",  x"28",  x"cd",  x"06",  x"cf",  x"e5",  x"eb", -- 70D0
         x"2b",  x"56",  x"2b",  x"5e",  x"e1",  x"cd",  x"29",  x"cd", -- 70D8
         x"cd",  x"db",  x"c8",  x"cd",  x"cc",  x"c8",  x"b4",  x"44", -- 70E0
         x"4d",  x"e3",  x"71",  x"23",  x"70",  x"c3",  x"84",  x"d1", -- 70E8
         x"cd",  x"45",  x"d1",  x"d5",  x"cd",  x"e1",  x"cd",  x"cd", -- 70F0
         x"29",  x"cd",  x"e3",  x"5e",  x"23",  x"56",  x"23",  x"7a", -- 70F8
         x"b3",  x"ca",  x"54",  x"c3",  x"7e",  x"23",  x"66",  x"6f", -- 7100
         x"e5",  x"2a",  x"df",  x"03",  x"e3",  x"22",  x"df",  x"03", -- 7108
         x"2a",  x"e3",  x"03",  x"e5",  x"2a",  x"e1",  x"03",  x"e5", -- 7110
         x"21",  x"e1",  x"03",  x"d5",  x"cd",  x"f7",  x"d6",  x"e1", -- 7118
         x"cd",  x"26",  x"cd",  x"cd",  x"be",  x"c8",  x"c2",  x"48", -- 7120
         x"c3",  x"e1",  x"22",  x"e1",  x"03",  x"e1",  x"22",  x"e3", -- 7128
         x"03",  x"e1",  x"22",  x"df",  x"03",  x"e1",  x"c9",  x"e5", -- 7130
         x"2a",  x"58",  x"03",  x"23",  x"7c",  x"b5",  x"e1",  x"c0", -- 7138
         x"1e",  x"16",  x"c3",  x"56",  x"c3",  x"cd",  x"cc",  x"c8", -- 7140
         x"a7",  x"3e",  x"80",  x"32",  x"cc",  x"03",  x"b6",  x"47", -- 7148
         x"cd",  x"0b",  x"cf",  x"c3",  x"29",  x"cd",  x"cd",  x"29", -- 7150
         x"cd",  x"cd",  x"34",  x"d8",  x"cd",  x"8a",  x"d1",  x"cd", -- 7158
         x"fe",  x"d2",  x"01",  x"57",  x"d3",  x"c5",  x"7e",  x"23", -- 7160
         x"23",  x"e5",  x"cd",  x"e1",  x"d1",  x"e1",  x"4e",  x"23", -- 7168
         x"46",  x"cd",  x"7e",  x"d1",  x"e5",  x"6f",  x"cd",  x"f2", -- 7170
         x"d2",  x"d1",  x"c9",  x"cd",  x"e1",  x"d1",  x"21",  x"c0", -- 7178
         x"03",  x"e5",  x"77",  x"23",  x"23",  x"73",  x"23",  x"72", -- 7180
         x"e1",  x"c9",  x"2b",  x"06",  x"22",  x"50",  x"e5",  x"0e", -- 7188
         x"ff",  x"23",  x"7e",  x"0c",  x"b7",  x"28",  x"06",  x"ba", -- 7190
         x"28",  x"03",  x"b8",  x"20",  x"f4",  x"fe",  x"22",  x"cc", -- 7198
         x"bd",  x"c8",  x"e3",  x"23",  x"eb",  x"79",  x"cd",  x"7e", -- 71A0
         x"d1",  x"11",  x"c0",  x"03",  x"2a",  x"b2",  x"03",  x"22", -- 71A8
         x"e5",  x"03",  x"3e",  x"01",  x"32",  x"ae",  x"03",  x"cd", -- 71B0
         x"fa",  x"d6",  x"cd",  x"89",  x"c6",  x"22",  x"b2",  x"03", -- 71B8
         x"e1",  x"7e",  x"c0",  x"1e",  x"1e",  x"c3",  x"56",  x"c3", -- 71C0
         x"23",  x"cd",  x"8a",  x"d1",  x"cd",  x"fe",  x"d2",  x"cd", -- 71C8
         x"ee",  x"d6",  x"1c",  x"1d",  x"c8",  x"0a",  x"cd",  x"ae", -- 71D0
         x"c6",  x"fe",  x"0d",  x"cc",  x"66",  x"cb",  x"03",  x"18", -- 71D8
         x"f2",  x"b7",  x"0e",  x"f1",  x"f5",  x"ed",  x"5b",  x"56", -- 71E0
         x"03",  x"2a",  x"c4",  x"03",  x"2f",  x"4f",  x"06",  x"ff", -- 71E8
         x"09",  x"23",  x"cd",  x"89",  x"c6",  x"38",  x"07",  x"22", -- 71F0
         x"c4",  x"03",  x"23",  x"eb",  x"f1",  x"c9",  x"f1",  x"1e", -- 71F8
         x"1a",  x"28",  x"c2",  x"bf",  x"f5",  x"01",  x"e3",  x"d1", -- 7200
         x"c5",  x"2a",  x"b0",  x"03",  x"22",  x"c4",  x"03",  x"21", -- 7208
         x"00",  x"00",  x"e5",  x"2a",  x"56",  x"03",  x"e5",  x"21", -- 7210
         x"b4",  x"03",  x"ed",  x"5b",  x"b2",  x"03",  x"cd",  x"89", -- 7218
         x"c6",  x"01",  x"1a",  x"d2",  x"20",  x"3f",  x"2a",  x"d7", -- 7220
         x"03",  x"ed",  x"5b",  x"d9",  x"03",  x"cd",  x"89",  x"c6", -- 7228
         x"28",  x"0a",  x"7e",  x"23",  x"23",  x"b7",  x"cd",  x"68", -- 7230
         x"d2",  x"18",  x"ee",  x"c1",  x"ed",  x"5b",  x"db",  x"03", -- 7238
         x"cd",  x"89",  x"c6",  x"28",  x"49",  x"cd",  x"ee",  x"d6", -- 7240
         x"7b",  x"e5",  x"09",  x"b7",  x"f2",  x"3b",  x"d2",  x"22", -- 7248
         x"c6",  x"03",  x"e1",  x"4e",  x"06",  x"00",  x"09",  x"09", -- 7250
         x"23",  x"ed",  x"5b",  x"c6",  x"03",  x"cd",  x"89",  x"c6", -- 7258
         x"28",  x"da",  x"01",  x"59",  x"d2",  x"c5",  x"f6",  x"80", -- 7260
         x"7e",  x"23",  x"23",  x"5e",  x"23",  x"56",  x"23",  x"f0", -- 7268
         x"b7",  x"c8",  x"44",  x"4d",  x"2a",  x"c4",  x"03",  x"cd", -- 7270
         x"89",  x"c6",  x"60",  x"69",  x"d8",  x"e1",  x"e3",  x"cd", -- 7278
         x"89",  x"c6",  x"e3",  x"e5",  x"60",  x"69",  x"d0",  x"c1", -- 7280
         x"f1",  x"f1",  x"e5",  x"d5",  x"c5",  x"c9",  x"d1",  x"e1", -- 7288
         x"7d",  x"b4",  x"c8",  x"2b",  x"46",  x"2b",  x"4e",  x"e5", -- 7290
         x"2b",  x"2b",  x"6e",  x"26",  x"00",  x"09",  x"50",  x"59", -- 7298
         x"2b",  x"44",  x"4d",  x"2a",  x"c4",  x"03",  x"cd",  x"ae", -- 72A0
         x"c4",  x"e1",  x"71",  x"23",  x"70",  x"69",  x"60",  x"2b", -- 72A8
         x"c3",  x"0c",  x"d2",  x"c5",  x"e5",  x"2a",  x"e5",  x"03", -- 72B0
         x"e3",  x"cd",  x"ad",  x"cd",  x"e3",  x"cd",  x"2a",  x"cd", -- 72B8
         x"7e",  x"e5",  x"2a",  x"e5",  x"03",  x"e5",  x"86",  x"1e", -- 72C0
         x"1c",  x"da",  x"56",  x"c3",  x"cd",  x"7b",  x"d1",  x"d1", -- 72C8
         x"cd",  x"02",  x"d3",  x"e3",  x"cd",  x"01",  x"d3",  x"e5", -- 72D0
         x"2a",  x"c2",  x"03",  x"eb",  x"cd",  x"e9",  x"d2",  x"cd", -- 72D8
         x"e9",  x"d2",  x"21",  x"46",  x"cd",  x"e3",  x"e5",  x"18", -- 72E0
         x"6f",  x"e1",  x"e3",  x"7e",  x"23",  x"23",  x"4e",  x"23", -- 72E8
         x"46",  x"6f",  x"2c",  x"2d",  x"c8",  x"0a",  x"12",  x"03", -- 72F0
         x"13",  x"18",  x"f8",  x"cd",  x"2a",  x"cd",  x"2a",  x"e5", -- 72F8
         x"03",  x"eb",  x"cd",  x"1b",  x"d3",  x"eb",  x"c0",  x"d5", -- 7300
         x"50",  x"59",  x"1b",  x"4e",  x"2a",  x"c4",  x"03",  x"cd", -- 7308
         x"89",  x"c6",  x"20",  x"05",  x"47",  x"09",  x"22",  x"c4", -- 7310
         x"03",  x"e1",  x"c9",  x"2a",  x"b2",  x"03",  x"2b",  x"46", -- 7318
         x"2b",  x"4e",  x"2b",  x"2b",  x"cd",  x"89",  x"c6",  x"c0", -- 7320
         x"22",  x"b2",  x"03",  x"c9",  x"01",  x"c0",  x"d0",  x"c5", -- 7328
         x"cd",  x"fb",  x"d2",  x"af",  x"57",  x"32",  x"ae",  x"03", -- 7330
         x"7e",  x"b7",  x"c9",  x"01",  x"c0",  x"d0",  x"c5",  x"cd", -- 7338
         x"30",  x"d3",  x"28",  x"55",  x"23",  x"23",  x"5e",  x"23", -- 7340
         x"56",  x"1a",  x"c9",  x"3e",  x"01",  x"cd",  x"7b",  x"d1", -- 7348
         x"cd",  x"24",  x"d4",  x"2a",  x"c2",  x"03",  x"73",  x"c1", -- 7350
         x"c3",  x"a9",  x"d1",  x"cd",  x"da",  x"d3",  x"af",  x"e3", -- 7358
         x"4f",  x"e5",  x"7e",  x"b8",  x"38",  x"02",  x"78",  x"11", -- 7360
         x"0e",  x"00",  x"c5",  x"cd",  x"e1",  x"d1",  x"c1",  x"e1", -- 7368
         x"e5",  x"23",  x"23",  x"46",  x"23",  x"66",  x"68",  x"06", -- 7370
         x"00",  x"09",  x"44",  x"4d",  x"cd",  x"7e",  x"d1",  x"6f", -- 7378
         x"cd",  x"f2",  x"d2",  x"d1",  x"cd",  x"02",  x"d3",  x"18", -- 7380
         x"cf",  x"cd",  x"da",  x"d3",  x"d1",  x"d5",  x"1a",  x"90", -- 7388
         x"18",  x"cd",  x"eb",  x"7e",  x"cd",  x"de",  x"d3",  x"04", -- 7390
         x"05",  x"ca",  x"67",  x"c9",  x"c5",  x"1e",  x"ff",  x"fe", -- 7398
         x"29",  x"28",  x"06",  x"cd",  x"d6",  x"c8",  x"cd",  x"21", -- 73A0
         x"d4",  x"cd",  x"db",  x"c8",  x"f1",  x"e3",  x"01",  x"61", -- 73A8
         x"d3",  x"c5",  x"3d",  x"be",  x"06",  x"00",  x"d0",  x"4f", -- 73B0
         x"7e",  x"91",  x"bb",  x"47",  x"d8",  x"43",  x"c9",  x"cd", -- 73B8
         x"30",  x"d3",  x"ca",  x"cf",  x"d4",  x"5f",  x"23",  x"23", -- 73C0
         x"7e",  x"23",  x"66",  x"6f",  x"e5",  x"19",  x"46",  x"72", -- 73C8
         x"e3",  x"c5",  x"7e",  x"cd",  x"a1",  x"d7",  x"c1",  x"e1", -- 73D0
         x"70",  x"c9",  x"eb",  x"cd",  x"db",  x"c8",  x"c1",  x"d1", -- 73D8
         x"c5",  x"43",  x"c9",  x"cd",  x"24",  x"d4",  x"4f",  x"ed", -- 73E0
         x"78",  x"c3",  x"c0",  x"d0",  x"cd",  x"14",  x"d4",  x"3a", -- 73E8
         x"06",  x"03",  x"4f",  x"7b",  x"ed",  x"79",  x"c9",  x"cd", -- 73F0
         x"14",  x"d4",  x"f5",  x"1e",  x"00",  x"cd",  x"be",  x"c8", -- 73F8
         x"28",  x"06",  x"cd",  x"d6",  x"c8",  x"cd",  x"21",  x"d4", -- 7400
         x"c1",  x"3a",  x"06",  x"03",  x"4f",  x"ed",  x"78",  x"ab", -- 7408
         x"a0",  x"28",  x"fa",  x"c9",  x"cd",  x"21",  x"d4",  x"32", -- 7410
         x"06",  x"03",  x"cd",  x"d6",  x"c8",  x"2b",  x"cd",  x"bd", -- 7418
         x"c8",  x"cd",  x"26",  x"cd",  x"cd",  x"61",  x"c9",  x"7a", -- 7420
         x"b7",  x"c2",  x"67",  x"c9",  x"cd",  x"be",  x"c8",  x"7b", -- 7428
         x"c9",  x"cd",  x"6f",  x"c9",  x"1a",  x"18",  x"b2",  x"cd", -- 7430
         x"6c",  x"c9",  x"d5",  x"cd",  x"d6",  x"c8",  x"cd",  x"21", -- 7438
         x"d4",  x"d1",  x"12",  x"c9",  x"cd",  x"6f",  x"c9",  x"eb", -- 7440
         x"46",  x"23",  x"7e",  x"c3",  x"b1",  x"d0",  x"cd",  x"6c", -- 7448
         x"c9",  x"d5",  x"cd",  x"d6",  x"c8",  x"cd",  x"6c",  x"c9", -- 7450
         x"e3",  x"73",  x"23",  x"72",  x"e1",  x"c9",  x"21",  x"04", -- 7458
         x"d9",  x"cd",  x"ee",  x"d6",  x"18",  x"09",  x"cd",  x"ee", -- 7460
         x"d6",  x"21",  x"c1",  x"d1",  x"cd",  x"c0",  x"d6",  x"78", -- 7468
         x"b7",  x"c8",  x"3a",  x"e8",  x"03",  x"b7",  x"ca",  x"e0", -- 7470
         x"d6",  x"90",  x"30",  x"0c",  x"2f",  x"3c",  x"eb",  x"cd", -- 7478
         x"c8",  x"d6",  x"eb",  x"cd",  x"e0",  x"d6",  x"c1",  x"d1", -- 7480
         x"fe",  x"19",  x"d0",  x"f5",  x"cd",  x"03",  x"d7",  x"67", -- 7488
         x"f1",  x"cd",  x"2a",  x"d5",  x"b4",  x"21",  x"e5",  x"03", -- 7490
         x"f2",  x"ab",  x"d4",  x"cd",  x"0a",  x"d5",  x"30",  x"4b", -- 7498
         x"23",  x"34",  x"28",  x"63",  x"2e",  x"01",  x"cd",  x"3e", -- 74A0
         x"d5",  x"18",  x"40",  x"af",  x"90",  x"47",  x"7e",  x"9b", -- 74A8
         x"5f",  x"23",  x"7e",  x"9a",  x"57",  x"23",  x"7e",  x"99", -- 74B0
         x"4f",  x"dc",  x"16",  x"d5",  x"68",  x"63",  x"af",  x"47", -- 74B8
         x"79",  x"b7",  x"20",  x"16",  x"4a",  x"54",  x"65",  x"6f", -- 74C0
         x"78",  x"d6",  x"08",  x"fe",  x"e0",  x"20",  x"f0",  x"af", -- 74C8
         x"32",  x"e8",  x"03",  x"c9",  x"05",  x"29",  x"cb",  x"12", -- 74D0
         x"cb",  x"11",  x"f2",  x"d4",  x"d4",  x"78",  x"5c",  x"45", -- 74D8
         x"b7",  x"28",  x"08",  x"21",  x"e8",  x"03",  x"86",  x"77", -- 74E0
         x"30",  x"e5",  x"c8",  x"78",  x"21",  x"e8",  x"03",  x"b7", -- 74E8
         x"fc",  x"fd",  x"d4",  x"46",  x"23",  x"7e",  x"e6",  x"80", -- 74F0
         x"a9",  x"4f",  x"c3",  x"e0",  x"d6",  x"1c",  x"c0",  x"14", -- 74F8
         x"c0",  x"0c",  x"c0",  x"0e",  x"80",  x"34",  x"c0",  x"c3", -- 7500
         x"53",  x"d6",  x"7e",  x"83",  x"5f",  x"23",  x"7e",  x"8a", -- 7508
         x"57",  x"23",  x"7e",  x"89",  x"4f",  x"c9",  x"21",  x"e9", -- 7510
         x"03",  x"7e",  x"2f",  x"77",  x"af",  x"6f",  x"90",  x"47", -- 7518
         x"7d",  x"9b",  x"5f",  x"7d",  x"9a",  x"57",  x"7d",  x"99", -- 7520
         x"4f",  x"c9",  x"06",  x"00",  x"d6",  x"08",  x"38",  x"07", -- 7528
         x"43",  x"5a",  x"51",  x"0e",  x"00",  x"18",  x"f5",  x"c6", -- 7530
         x"09",  x"6f",  x"af",  x"2d",  x"c8",  x"79",  x"1f",  x"4f", -- 7538
         x"cb",  x"1a",  x"cb",  x"1b",  x"cb",  x"18",  x"18",  x"f2", -- 7540
         x"00",  x"00",  x"00",  x"81",  x"03",  x"aa",  x"56",  x"19", -- 7548
         x"80",  x"f1",  x"22",  x"76",  x"80",  x"45",  x"aa",  x"38", -- 7550
         x"82",  x"cd",  x"97",  x"d6",  x"b7",  x"ea",  x"67",  x"c9", -- 7558
         x"21",  x"e8",  x"03",  x"7e",  x"01",  x"35",  x"80",  x"11", -- 7560
         x"f3",  x"04",  x"90",  x"f5",  x"70",  x"d5",  x"c5",  x"cd", -- 7568
         x"6f",  x"d4",  x"c1",  x"d1",  x"04",  x"cd",  x"f5",  x"d5", -- 7570
         x"21",  x"48",  x"d5",  x"cd",  x"66",  x"d4",  x"21",  x"4c", -- 7578
         x"d5",  x"cd",  x"ce",  x"d9",  x"01",  x"80",  x"80",  x"11", -- 7580
         x"00",  x"00",  x"cd",  x"6f",  x"d4",  x"f1",  x"cd",  x"0b", -- 7588
         x"d8",  x"01",  x"31",  x"80",  x"11",  x"18",  x"72",  x"21", -- 7590
         x"c1",  x"d1",  x"cd",  x"97",  x"d6",  x"c8",  x"2e",  x"00", -- 7598
         x"cd",  x"58",  x"d6",  x"79",  x"32",  x"f7",  x"03",  x"eb", -- 75A0
         x"22",  x"f8",  x"03",  x"01",  x"00",  x"00",  x"50",  x"58", -- 75A8
         x"21",  x"bc",  x"d4",  x"e5",  x"21",  x"bc",  x"d5",  x"e5", -- 75B0
         x"e5",  x"21",  x"e5",  x"03",  x"7e",  x"23",  x"b7",  x"28", -- 75B8
         x"21",  x"e5",  x"2e",  x"08",  x"1f",  x"67",  x"79",  x"30", -- 75C0
         x"0b",  x"e5",  x"2a",  x"f8",  x"03",  x"19",  x"eb",  x"e1", -- 75C8
         x"3a",  x"f7",  x"03",  x"89",  x"1f",  x"4f",  x"cb",  x"1a", -- 75D0
         x"cb",  x"1b",  x"cb",  x"18",  x"2d",  x"7c",  x"20",  x"e4", -- 75D8
         x"e1",  x"c9",  x"43",  x"5a",  x"51",  x"4f",  x"c9",  x"cd", -- 75E0
         x"c8",  x"d6",  x"01",  x"20",  x"84",  x"11",  x"00",  x"00", -- 75E8
         x"cd",  x"e0",  x"d6",  x"c1",  x"d1",  x"cd",  x"97",  x"d6", -- 75F0
         x"ca",  x"4b",  x"c3",  x"2e",  x"ff",  x"cd",  x"58",  x"d6", -- 75F8
         x"34",  x"34",  x"2b",  x"7e",  x"32",  x"14",  x"03",  x"2b", -- 7600
         x"7e",  x"32",  x"10",  x"03",  x"2b",  x"7e",  x"32",  x"0c", -- 7608
         x"03",  x"41",  x"eb",  x"af",  x"4f",  x"57",  x"5f",  x"32", -- 7610
         x"17",  x"03",  x"e5",  x"c5",  x"7d",  x"cd",  x"0b",  x"03", -- 7618
         x"de",  x"00",  x"3f",  x"30",  x"07",  x"32",  x"17",  x"03", -- 7620
         x"f1",  x"f1",  x"37",  x"d2",  x"c1",  x"e1",  x"79",  x"3c", -- 7628
         x"3d",  x"1f",  x"fa",  x"ec",  x"d4",  x"17",  x"cb",  x"13", -- 7630
         x"cb",  x"12",  x"cb",  x"11",  x"29",  x"cb",  x"10",  x"3a", -- 7638
         x"17",  x"03",  x"17",  x"32",  x"17",  x"03",  x"79",  x"b2", -- 7640
         x"b3",  x"20",  x"cf",  x"e5",  x"21",  x"e8",  x"03",  x"35", -- 7648
         x"e1",  x"20",  x"c7",  x"1e",  x"0a",  x"c3",  x"56",  x"c3", -- 7650
         x"78",  x"b7",  x"ca",  x"7c",  x"d6",  x"7d",  x"21",  x"e8", -- 7658
         x"03",  x"ae",  x"80",  x"47",  x"1f",  x"a8",  x"78",  x"f2", -- 7660
         x"7b",  x"d6",  x"c6",  x"80",  x"77",  x"ca",  x"e0",  x"d5", -- 7668
         x"cd",  x"03",  x"d7",  x"77",  x"2b",  x"c9",  x"cd",  x"97", -- 7670
         x"d6",  x"2f",  x"e1",  x"b7",  x"e1",  x"f2",  x"cf",  x"d4", -- 7678
         x"18",  x"d1",  x"cd",  x"eb",  x"d6",  x"78",  x"b7",  x"c8", -- 7680
         x"c6",  x"02",  x"38",  x"c7",  x"47",  x"cd",  x"6f",  x"d4", -- 7688
         x"21",  x"e8",  x"03",  x"34",  x"c0",  x"18",  x"bc",  x"3a", -- 7690
         x"e8",  x"03",  x"b7",  x"c8",  x"3a",  x"e7",  x"03",  x"fe", -- 7698
         x"2f",  x"17",  x"9f",  x"c0",  x"3c",  x"c9",  x"cd",  x"97", -- 76A0
         x"d6",  x"06",  x"88",  x"11",  x"00",  x"00",  x"21",  x"e8", -- 76A8
         x"03",  x"4f",  x"70",  x"06",  x"00",  x"23",  x"36",  x"80", -- 76B0
         x"17",  x"c3",  x"b9",  x"d4",  x"cd",  x"97",  x"d6",  x"f0", -- 76B8
         x"21",  x"e7",  x"03",  x"7e",  x"ee",  x"80",  x"77",  x"c9", -- 76C0
         x"eb",  x"2a",  x"e5",  x"03",  x"e3",  x"e5",  x"2a",  x"e7", -- 76C8
         x"03",  x"e3",  x"e5",  x"eb",  x"c9",  x"01",  x"49",  x"82", -- 76D0
         x"11",  x"db",  x"0f",  x"18",  x"03",  x"cd",  x"ee",  x"d6", -- 76D8
         x"ed",  x"53",  x"e5",  x"03",  x"ed",  x"43",  x"e7",  x"03", -- 76E0
         x"50",  x"59",  x"c9",  x"21",  x"e5",  x"03",  x"5e",  x"23", -- 76E8
         x"56",  x"23",  x"4e",  x"23",  x"46",  x"23",  x"c9",  x"11", -- 76F0
         x"e5",  x"03",  x"06",  x"04",  x"1a",  x"77",  x"13",  x"23", -- 76F8
         x"10",  x"fa",  x"c9",  x"21",  x"e7",  x"03",  x"7e",  x"07", -- 7700
         x"37",  x"1f",  x"77",  x"3f",  x"1f",  x"23",  x"23",  x"77", -- 7708
         x"79",  x"07",  x"37",  x"1f",  x"4f",  x"1f",  x"ae",  x"c9", -- 7710
         x"78",  x"b7",  x"ca",  x"97",  x"d6",  x"21",  x"a0",  x"d6", -- 7718
         x"e5",  x"cd",  x"97",  x"d6",  x"79",  x"c8",  x"21",  x"e7", -- 7720
         x"03",  x"ae",  x"79",  x"f8",  x"cd",  x"32",  x"d7",  x"1f", -- 7728
         x"a9",  x"c9",  x"23",  x"78",  x"be",  x"c0",  x"2b",  x"79", -- 7730
         x"be",  x"c0",  x"2b",  x"7a",  x"be",  x"c0",  x"2b",  x"7b", -- 7738
         x"96",  x"c0",  x"e1",  x"e1",  x"c9",  x"47",  x"4f",  x"57", -- 7740
         x"5f",  x"b7",  x"c8",  x"e5",  x"cd",  x"eb",  x"d6",  x"cd", -- 7748
         x"03",  x"d7",  x"ae",  x"67",  x"fc",  x"69",  x"d7",  x"3e", -- 7750
         x"98",  x"90",  x"cd",  x"2a",  x"d5",  x"7c",  x"17",  x"dc", -- 7758
         x"fd",  x"d4",  x"06",  x"00",  x"dc",  x"16",  x"d5",  x"e1", -- 7760
         x"c9",  x"1b",  x"7a",  x"a3",  x"3c",  x"c0",  x"0b",  x"c9", -- 7768
         x"21",  x"e8",  x"03",  x"7e",  x"fe",  x"98",  x"3a",  x"e5", -- 7770
         x"03",  x"d0",  x"7e",  x"cd",  x"45",  x"d7",  x"36",  x"98", -- 7778
         x"7b",  x"f5",  x"79",  x"17",  x"cd",  x"b9",  x"d4",  x"f1", -- 7780
         x"c9",  x"21",  x"00",  x"00",  x"78",  x"b1",  x"c8",  x"3e", -- 7788
         x"10",  x"29",  x"38",  x"06",  x"eb",  x"29",  x"eb",  x"30", -- 7790
         x"04",  x"09",  x"da",  x"0b",  x"d0",  x"3d",  x"20",  x"f1", -- 7798
         x"c9",  x"fe",  x"2d",  x"f5",  x"28",  x"05",  x"fe",  x"2b", -- 77A0
         x"28",  x"01",  x"2b",  x"cd",  x"cf",  x"d4",  x"47",  x"57", -- 77A8
         x"5f",  x"2f",  x"4f",  x"cd",  x"bd",  x"c8",  x"38",  x"3d", -- 77B0
         x"fe",  x"2e",  x"28",  x"16",  x"fe",  x"45",  x"20",  x"15", -- 77B8
         x"cd",  x"bd",  x"c8",  x"cd",  x"4d",  x"ce",  x"cd",  x"bd", -- 77C0
         x"c8",  x"38",  x"4b",  x"14",  x"20",  x"07",  x"af",  x"93", -- 77C8
         x"5f",  x"0c",  x"0c",  x"28",  x"de",  x"e5",  x"7b",  x"90", -- 77D0
         x"f4",  x"ed",  x"d7",  x"f2",  x"e4",  x"d7",  x"f5",  x"cd", -- 77D8
         x"e7",  x"d5",  x"f1",  x"3c",  x"20",  x"f2",  x"d1",  x"f1", -- 77E0
         x"cc",  x"c0",  x"d6",  x"eb",  x"c9",  x"c8",  x"f5",  x"cd", -- 77E8
         x"82",  x"d6",  x"f1",  x"3d",  x"c9",  x"d5",  x"57",  x"78", -- 77F0
         x"89",  x"47",  x"c5",  x"e5",  x"d5",  x"cd",  x"82",  x"d6", -- 77F8
         x"f1",  x"d6",  x"30",  x"cd",  x"0b",  x"d8",  x"e1",  x"c1", -- 7800
         x"d1",  x"18",  x"a8",  x"cd",  x"c8",  x"d6",  x"cd",  x"a9", -- 7808
         x"d6",  x"c1",  x"d1",  x"c3",  x"6f",  x"d4",  x"7b",  x"07", -- 7810
         x"07",  x"83",  x"07",  x"86",  x"d6",  x"30",  x"5f",  x"18", -- 7818
         x"a5",  x"e5",  x"21",  x"0d",  x"c3",  x"cd",  x"c9",  x"d1", -- 7820
         x"e1",  x"eb",  x"af",  x"06",  x"98",  x"cd",  x"ae",  x"d6", -- 7828
         x"21",  x"c8",  x"d1",  x"e5",  x"21",  x"ea",  x"03",  x"e5", -- 7830
         x"cd",  x"97",  x"d6",  x"36",  x"20",  x"f2",  x"42",  x"d8", -- 7838
         x"36",  x"2d",  x"23",  x"36",  x"30",  x"ca",  x"ef",  x"d8", -- 7840
         x"e5",  x"fc",  x"c0",  x"d6",  x"af",  x"f5",  x"cd",  x"f5", -- 7848
         x"d8",  x"01",  x"43",  x"91",  x"11",  x"f8",  x"4f",  x"cd", -- 7850
         x"18",  x"d7",  x"b7",  x"e2",  x"6e",  x"d8",  x"f1",  x"cd", -- 7858
         x"ee",  x"d7",  x"f5",  x"18",  x"ec",  x"cd",  x"e7",  x"d5", -- 7860
         x"f1",  x"3c",  x"f5",  x"cd",  x"f5",  x"d8",  x"cd",  x"5e", -- 7868
         x"d4",  x"3c",  x"cd",  x"45",  x"d7",  x"cd",  x"e0",  x"d6", -- 7870
         x"01",  x"06",  x"03",  x"f1",  x"81",  x"3c",  x"fa",  x"89", -- 7878
         x"d8",  x"fe",  x"08",  x"30",  x"04",  x"3c",  x"47",  x"3e", -- 7880
         x"02",  x"3d",  x"3d",  x"e1",  x"f5",  x"11",  x"08",  x"d9", -- 7888
         x"05",  x"20",  x"06",  x"36",  x"2e",  x"23",  x"36",  x"30", -- 7890
         x"23",  x"05",  x"36",  x"2e",  x"cc",  x"f5",  x"d6",  x"c5", -- 7898
         x"e5",  x"d5",  x"cd",  x"eb",  x"d6",  x"e1",  x"06",  x"2f", -- 78A0
         x"04",  x"7b",  x"96",  x"5f",  x"23",  x"7a",  x"9e",  x"57", -- 78A8
         x"23",  x"79",  x"9e",  x"4f",  x"2b",  x"2b",  x"30",  x"f0", -- 78B0
         x"cd",  x"0a",  x"d5",  x"23",  x"cd",  x"e0",  x"d6",  x"eb", -- 78B8
         x"e1",  x"70",  x"23",  x"c1",  x"0d",  x"20",  x"d2",  x"05", -- 78C0
         x"28",  x"0b",  x"2b",  x"7e",  x"fe",  x"30",  x"28",  x"fa", -- 78C8
         x"fe",  x"2e",  x"c4",  x"f5",  x"d6",  x"f1",  x"28",  x"1a", -- 78D0
         x"36",  x"45",  x"23",  x"36",  x"2b",  x"f2",  x"e4",  x"d8", -- 78D8
         x"36",  x"2d",  x"2f",  x"3c",  x"06",  x"2f",  x"04",  x"d6", -- 78E0
         x"0a",  x"30",  x"fb",  x"c6",  x"3a",  x"23",  x"70",  x"23", -- 78E8
         x"77",  x"23",  x"71",  x"e1",  x"c9",  x"01",  x"74",  x"94", -- 78F0
         x"11",  x"f7",  x"23",  x"cd",  x"18",  x"d7",  x"b7",  x"e1", -- 78F8
         x"e2",  x"65",  x"d8",  x"e9",  x"00",  x"00",  x"00",  x"80", -- 7900
         x"a0",  x"86",  x"01",  x"10",  x"27",  x"00",  x"e8",  x"03", -- 7908
         x"00",  x"64",  x"00",  x"00",  x"0a",  x"00",  x"00",  x"01", -- 7910
         x"00",  x"00",  x"21",  x"c0",  x"d6",  x"e3",  x"e9",  x"cd", -- 7918
         x"c8",  x"d6",  x"21",  x"04",  x"d9",  x"cd",  x"dd",  x"d6", -- 7920
         x"c1",  x"d1",  x"cd",  x"97",  x"d6",  x"78",  x"ca",  x"6d", -- 7928
         x"d9",  x"f2",  x"38",  x"d9",  x"b7",  x"ca",  x"4b",  x"c3", -- 7930
         x"b7",  x"ca",  x"d0",  x"d4",  x"d5",  x"c5",  x"79",  x"f6", -- 7938
         x"7f",  x"cd",  x"eb",  x"d6",  x"f2",  x"55",  x"d9",  x"d5", -- 7940
         x"c5",  x"cd",  x"70",  x"d7",  x"c1",  x"d1",  x"f5",  x"cd", -- 7948
         x"18",  x"d7",  x"e1",  x"7c",  x"1f",  x"e1",  x"22",  x"e7", -- 7950
         x"03",  x"e1",  x"22",  x"e5",  x"03",  x"dc",  x"1a",  x"d9", -- 7958
         x"cc",  x"c0",  x"d6",  x"d5",  x"c5",  x"cd",  x"59",  x"d5", -- 7960
         x"c1",  x"d1",  x"cd",  x"9a",  x"d5",  x"cd",  x"c8",  x"d6", -- 7968
         x"01",  x"38",  x"81",  x"11",  x"3b",  x"aa",  x"cd",  x"9a", -- 7970
         x"d5",  x"3a",  x"e8",  x"03",  x"fe",  x"88",  x"d2",  x"76", -- 7978
         x"d6",  x"cd",  x"70",  x"d7",  x"c6",  x"80",  x"c6",  x"02", -- 7980
         x"da",  x"76",  x"d6",  x"f5",  x"21",  x"48",  x"d5",  x"cd", -- 7988
         x"61",  x"d4",  x"cd",  x"91",  x"d5",  x"f1",  x"c1",  x"d1", -- 7990
         x"f5",  x"cd",  x"6c",  x"d4",  x"cd",  x"c0",  x"d6",  x"21", -- 7998
         x"ad",  x"d9",  x"cd",  x"dd",  x"d9",  x"11",  x"00",  x"00", -- 79A0
         x"c1",  x"4a",  x"c3",  x"9a",  x"d5",  x"08",  x"40",  x"2e", -- 79A8
         x"94",  x"74",  x"70",  x"4f",  x"2e",  x"77",  x"6e",  x"02", -- 79B0
         x"88",  x"7a",  x"e6",  x"a0",  x"2a",  x"7c",  x"50",  x"aa", -- 79B8
         x"aa",  x"7e",  x"ff",  x"ff",  x"7f",  x"7f",  x"00",  x"00", -- 79C0
         x"80",  x"81",  x"00",  x"00",  x"00",  x"81",  x"cd",  x"c8", -- 79C8
         x"d6",  x"11",  x"98",  x"d5",  x"d5",  x"e5",  x"cd",  x"eb", -- 79D0
         x"d6",  x"cd",  x"9a",  x"d5",  x"e1",  x"cd",  x"c8",  x"d6", -- 79D8
         x"7e",  x"23",  x"cd",  x"dd",  x"d6",  x"06",  x"f1",  x"c1", -- 79E0
         x"d1",  x"3d",  x"c8",  x"d5",  x"c5",  x"f5",  x"e5",  x"cd", -- 79E8
         x"9a",  x"d5",  x"e1",  x"cd",  x"ee",  x"d6",  x"e5",  x"cd", -- 79F0
         x"6f",  x"d4",  x"e1",  x"18",  x"e9",  x"cd",  x"97",  x"d6", -- 79F8
         x"21",  x"1b",  x"03",  x"fa",  x"5d",  x"da",  x"21",  x"3c", -- 7A00
         x"03",  x"cd",  x"dd",  x"d6",  x"21",  x"1b",  x"03",  x"c8", -- 7A08
         x"86",  x"e6",  x"07",  x"06",  x"00",  x"77",  x"23",  x"87", -- 7A10
         x"87",  x"4f",  x"09",  x"cd",  x"ee",  x"d6",  x"cd",  x"9a", -- 7A18
         x"d5",  x"3a",  x"1a",  x"03",  x"3c",  x"e6",  x"03",  x"06", -- 7A20
         x"00",  x"fe",  x"01",  x"88",  x"32",  x"1a",  x"03",  x"21", -- 7A28
         x"60",  x"da",  x"87",  x"87",  x"4f",  x"09",  x"cd",  x"61", -- 7A30
         x"d4",  x"cd",  x"eb",  x"d6",  x"7b",  x"59",  x"ee",  x"4f", -- 7A38
         x"4f",  x"36",  x"80",  x"2b",  x"46",  x"36",  x"80",  x"21", -- 7A40
         x"19",  x"03",  x"34",  x"7e",  x"d6",  x"ab",  x"20",  x"04", -- 7A48
         x"77",  x"0c",  x"15",  x"1c",  x"cd",  x"bc",  x"d4",  x"21", -- 7A50
         x"3c",  x"03",  x"c3",  x"f7",  x"d6",  x"77",  x"2b",  x"77", -- 7A58
         x"2b",  x"77",  x"18",  x"d5",  x"68",  x"b1",  x"46",  x"68", -- 7A60
         x"99",  x"e9",  x"92",  x"69",  x"10",  x"d1",  x"75",  x"68", -- 7A68
         x"21",  x"ba",  x"da",  x"cd",  x"61",  x"d4",  x"cd",  x"c8", -- 7A70
         x"d6",  x"01",  x"49",  x"83",  x"11",  x"db",  x"0f",  x"cd", -- 7A78
         x"e0",  x"d6",  x"c1",  x"d1",  x"cd",  x"f5",  x"d5",  x"cd", -- 7A80
         x"c8",  x"d6",  x"cd",  x"70",  x"d7",  x"c1",  x"d1",  x"cd", -- 7A88
         x"6c",  x"d4",  x"21",  x"be",  x"da",  x"cd",  x"66",  x"d4", -- 7A90
         x"cd",  x"97",  x"d6",  x"37",  x"f2",  x"a6",  x"da",  x"cd", -- 7A98
         x"5e",  x"d4",  x"cd",  x"97",  x"d6",  x"b7",  x"f5",  x"f4", -- 7AA0
         x"c0",  x"d6",  x"21",  x"be",  x"da",  x"cd",  x"61",  x"d4", -- 7AA8
         x"f1",  x"d4",  x"c0",  x"d6",  x"21",  x"c2",  x"da",  x"c3", -- 7AB0
         x"ce",  x"d9",  x"db",  x"0f",  x"49",  x"81",  x"00",  x"00", -- 7AB8
         x"00",  x"7f",  x"05",  x"ba",  x"d7",  x"1e",  x"86",  x"64", -- 7AC0
         x"26",  x"99",  x"87",  x"58",  x"34",  x"23",  x"87",  x"e0", -- 7AC8
         x"5d",  x"a5",  x"86",  x"da",  x"0f",  x"49",  x"83",  x"cd", -- 7AD0
         x"c8",  x"d6",  x"cd",  x"76",  x"da",  x"c1",  x"e1",  x"cd", -- 7AD8
         x"c8",  x"d6",  x"eb",  x"cd",  x"e0",  x"d6",  x"cd",  x"70", -- 7AE0
         x"da",  x"c3",  x"f3",  x"d5",  x"cd",  x"97",  x"d6",  x"fc", -- 7AE8
         x"1a",  x"d9",  x"fc",  x"c0",  x"d6",  x"3a",  x"e8",  x"03", -- 7AF0
         x"fe",  x"81",  x"da",  x"09",  x"db",  x"01",  x"00",  x"81", -- 7AF8
         x"51",  x"59",  x"cd",  x"f5",  x"d5",  x"21",  x"66",  x"d4", -- 7B00
         x"e5",  x"21",  x"13",  x"db",  x"cd",  x"ce",  x"d9",  x"21", -- 7B08
         x"ba",  x"da",  x"c9",  x"09",  x"4a",  x"d7",  x"3b",  x"78", -- 7B10
         x"02",  x"6e",  x"84",  x"7b",  x"fe",  x"c1",  x"2f",  x"7c", -- 7B18
         x"74",  x"31",  x"9a",  x"7d",  x"84",  x"3d",  x"5a",  x"7d", -- 7B20
         x"c8",  x"7f",  x"91",  x"7e",  x"e4",  x"bb",  x"4c",  x"7e", -- 7B28
         x"6c",  x"aa",  x"aa",  x"7f",  x"00",  x"00",  x"00",  x"81", -- 7B30
         x"cd",  x"49",  x"db",  x"28",  x"03",  x"cd",  x"6c",  x"c9", -- 7B38
         x"e5",  x"21",  x"47",  x"db",  x"e5",  x"eb",  x"e9",  x"e1", -- 7B40
         x"c9",  x"fe",  x"ae",  x"c0",  x"11",  x"00",  x"00",  x"cd", -- 7B48
         x"bd",  x"c8",  x"c8",  x"38",  x"0b",  x"fe",  x"94",  x"28", -- 7B50
         x"16",  x"fe",  x"47",  x"d2",  x"48",  x"c3",  x"d6",  x"07", -- 7B58
         x"d6",  x"30",  x"da",  x"48",  x"c3",  x"eb",  x"29",  x"29", -- 7B60
         x"29",  x"29",  x"b5",  x"6f",  x"eb",  x"18",  x"e0",  x"7b", -- 7B68
         x"87",  x"87",  x"87",  x"87",  x"f6",  x"0d",  x"57",  x"1e", -- 7B70
         x"ef",  x"18",  x"d4",  x"d5",  x"e5",  x"36",  x"00",  x"23", -- 7B78
         x"cd",  x"89",  x"c6",  x"20",  x"f8",  x"e3",  x"e5",  x"cd", -- 7B80
         x"fe",  x"d2",  x"cd",  x"09",  x"d2",  x"2a",  x"c4",  x"03", -- 7B88
         x"ed",  x"5b",  x"56",  x"03",  x"af",  x"ed",  x"52",  x"d1", -- 7B90
         x"e3",  x"ed",  x"52",  x"e5",  x"cd",  x"28",  x"dd",  x"4f", -- 7B98
         x"cd",  x"e4",  x"dd",  x"47",  x"e1",  x"cd",  x"e4",  x"dd", -- 7BA0
         x"12",  x"13",  x"2b",  x"7d",  x"b4",  x"20",  x"f6",  x"e1", -- 7BA8
         x"cd",  x"e4",  x"dd",  x"5f",  x"cd",  x"e4",  x"dd",  x"57", -- 7BB0
         x"af",  x"ed",  x"52",  x"38",  x"44",  x"2a",  x"56",  x"03", -- 7BB8
         x"23",  x"cd",  x"e4",  x"dd",  x"77",  x"23",  x"1b",  x"7b", -- 7BC0
         x"b2",  x"20",  x"f6",  x"d1",  x"e3",  x"c5",  x"cd",  x"f8", -- 7BC8
         x"dc",  x"e3",  x"ed",  x"42",  x"20",  x"2d",  x"e1",  x"cd", -- 7BD0
         x"77",  x"dd",  x"e3",  x"2b",  x"d5",  x"ed",  x"5b",  x"c4", -- 7BD8
         x"03",  x"ed",  x"b8",  x"ed",  x"53",  x"c4",  x"03",  x"e1", -- 7BE0
         x"42",  x"4b",  x"03",  x"d1",  x"2b",  x"70",  x"2b",  x"71", -- 7BE8
         x"2b",  x"35",  x"03",  x"20",  x"fc",  x"0b",  x"2b",  x"cd", -- 7BF0
         x"89",  x"c6",  x"20",  x"f0",  x"e1",  x"cd",  x"fd",  x"dd", -- 7BF8
         x"c9",  x"d1",  x"e1",  x"36",  x"00",  x"23",  x"cd",  x"89", -- 7C00
         x"c6",  x"20",  x"f8",  x"18",  x"29",  x"cd",  x"87",  x"dc", -- 7C08
         x"e5",  x"e2",  x"7b",  x"db",  x"eb",  x"ed",  x"52",  x"e5", -- 7C10
         x"cd",  x"28",  x"dd",  x"4f",  x"cd",  x"e4",  x"dd",  x"47", -- 7C18
         x"e1",  x"cd",  x"e4",  x"dd",  x"12",  x"13",  x"2b",  x"7d", -- 7C20
         x"b4",  x"20",  x"f6",  x"e1",  x"c5",  x"cd",  x"f8",  x"dc", -- 7C28
         x"e1",  x"ed",  x"42",  x"e1",  x"28",  x"c7",  x"cd",  x"1d", -- 7C30
         x"de",  x"21",  x"3f",  x"dc",  x"c3",  x"71",  x"c3",  x"42", -- 7C38
         x"41",  x"44",  x"00",  x"fe",  x"ae",  x"28",  x"c6",  x"cd", -- 7C40
         x"b0",  x"dc",  x"ed",  x"5b",  x"d7",  x"03",  x"1b",  x"1b", -- 7C48
         x"21",  x"00",  x"00",  x"39",  x"01",  x"d1",  x"ff",  x"ed", -- 7C50
         x"52",  x"09",  x"44",  x"4d",  x"cd",  x"28",  x"dd",  x"6f", -- 7C58
         x"cd",  x"e4",  x"dd",  x"67",  x"e5",  x"ed",  x"42",  x"e1", -- 7C60
         x"d2",  x"3e",  x"c3",  x"cd",  x"e4",  x"dd",  x"12",  x"13", -- 7C68
         x"2b",  x"7d",  x"b4",  x"20",  x"f6",  x"ed",  x"53",  x"d7", -- 7C70
         x"03",  x"21",  x"12",  x"c3",  x"cd",  x"c9",  x"d1",  x"c3", -- 7C78
         x"8a",  x"c4",  x"1e",  x"26",  x"c3",  x"56",  x"c3",  x"cd", -- 7C80
         x"ac",  x"dc",  x"e1",  x"cd",  x"cc",  x"c8",  x"3b",  x"3e", -- 7C88
         x"01",  x"32",  x"cc",  x"03",  x"cd",  x"06",  x"cf",  x"32", -- 7C90
         x"cc",  x"03",  x"e3",  x"e5",  x"60",  x"69",  x"eb",  x"19", -- 7C98
         x"eb",  x"4e",  x"06",  x"00",  x"09",  x"09",  x"23",  x"3a", -- 7CA0
         x"ae",  x"03",  x"b7",  x"c9",  x"3e",  x"d4",  x"23",  x"01", -- 7CA8
         x"3e",  x"d3",  x"f5",  x"3a",  x"5d",  x"03",  x"a7",  x"3e", -- 7CB0
         x"00",  x"32",  x"5d",  x"03",  x"28",  x"04",  x"f1",  x"c6", -- 7CB8
         x"04",  x"f5",  x"cd",  x"be",  x"c8",  x"cd",  x"3a",  x"cd", -- 7CC0
         x"f1",  x"e3",  x"e5",  x"f5",  x"cd",  x"3f",  x"d3",  x"21", -- 7CC8
         x"f7",  x"03",  x"06",  x"0d",  x"2b",  x"36",  x"20",  x"10", -- 7CD0
         x"fb",  x"d5",  x"11",  x"82",  x"dc",  x"73",  x"23",  x"72", -- 7CD8
         x"d1",  x"23",  x"f1",  x"77",  x"23",  x"77",  x"23",  x"77", -- 7CE0
         x"23",  x"eb",  x"06",  x"00",  x"79",  x"fe",  x"09",  x"38", -- 7CE8
         x"04",  x"0d",  x"23",  x"18",  x"f7",  x"ed",  x"b0",  x"c9", -- 7CF0
         x"e5",  x"af",  x"47",  x"86",  x"cd",  x"03",  x"dd",  x"20", -- 7CF8
         x"fa",  x"e1",  x"c9",  x"4f",  x"30",  x"01",  x"04",  x"23", -- 7D00
         x"cd",  x"89",  x"c6",  x"79",  x"c9",  x"f5",  x"3a",  x"07", -- 7D08
         x"03",  x"cb",  x"4f",  x"cb",  x"cf",  x"32",  x"07",  x"03", -- 7D10
         x"3e",  x"13",  x"20",  x"02",  x"c6",  x"08",  x"32",  x"08", -- 7D18
         x"03",  x"21",  x"ea",  x"03",  x"f1",  x"c3",  x"d5",  x"dd", -- 7D20
         x"3a",  x"07",  x"03",  x"cb",  x"47",  x"cb",  x"c7",  x"32", -- 7D28
         x"07",  x"03",  x"3e",  x"12",  x"20",  x"02",  x"c6",  x"08", -- 7D30
         x"32",  x"09",  x"03",  x"21",  x"ea",  x"03",  x"c3",  x"e4", -- 7D38
         x"dd",  x"fe",  x"ae",  x"28",  x"24",  x"cd",  x"97",  x"c6", -- 7D40
         x"cd",  x"b0",  x"dc",  x"2a",  x"d7",  x"03",  x"11",  x"ff", -- 7D48
         x"fb",  x"19",  x"44",  x"4d",  x"11",  x"01",  x"04",  x"cd", -- 7D50
         x"b5",  x"dd",  x"e1",  x"e5",  x"21",  x"07",  x"03",  x"cb", -- 7D58
         x"8e",  x"11",  x"43",  x"03",  x"cd",  x"f6",  x"df",  x"e1", -- 7D60
         x"c9",  x"cd",  x"87",  x"dc",  x"e2",  x"89",  x"dd",  x"cd", -- 7D68
         x"f8",  x"dc",  x"eb",  x"ed",  x"52",  x"18",  x"e0",  x"e5", -- 7D70
         x"01",  x"00",  x"00",  x"7e",  x"23",  x"77",  x"34",  x"81", -- 7D78
         x"23",  x"23",  x"cd",  x"03",  x"dd",  x"20",  x"f4",  x"e1", -- 7D80
         x"c9",  x"cd",  x"77",  x"dd",  x"c5",  x"cd",  x"f8",  x"dc", -- 7D88
         x"eb",  x"ed",  x"52",  x"cd",  x"b5",  x"dd",  x"c1",  x"79", -- 7D90
         x"cd",  x"d5",  x"dd",  x"78",  x"eb",  x"cd",  x"d5",  x"dd", -- 7D98
         x"2b",  x"2b",  x"78",  x"b1",  x"28",  x"b4",  x"56",  x"2b", -- 7DA0
         x"5e",  x"2b",  x"35",  x"28",  x"f3",  x"1a",  x"cd",  x"d5", -- 7DA8
         x"dd",  x"13",  x"0b",  x"18",  x"f5",  x"23",  x"e5",  x"79", -- 7DB0
         x"cd",  x"0d",  x"dd",  x"78",  x"e1",  x"cd",  x"d5",  x"dd", -- 7DB8
         x"2b",  x"7d",  x"b4",  x"1a",  x"13",  x"20",  x"f6",  x"c9", -- 7DC0
         x"3a",  x"08",  x"03",  x"e6",  x"07",  x"d6",  x"01",  x"c9", -- 7DC8
         x"cd",  x"1d",  x"de",  x"3e",  x"0c",  x"f5",  x"d5",  x"57", -- 7DD0
         x"3a",  x"08",  x"03",  x"5f",  x"7a",  x"cd",  x"f6",  x"df", -- 7DD8
         x"7b",  x"d1",  x"18",  x"3c",  x"d5",  x"3a",  x"09",  x"03", -- 7DE0
         x"5f",  x"cd",  x"f6",  x"df",  x"7b",  x"32",  x"09",  x"03", -- 7DE8
         x"7a",  x"18",  x"06",  x"d5",  x"1e",  x"80",  x"cd",  x"f6", -- 7DF0
         x"df",  x"cb",  x"7b",  x"d1",  x"c9",  x"f5",  x"e5",  x"d5", -- 7DF8
         x"c5",  x"11",  x"42",  x"03",  x"06",  x"06",  x"7a",  x"21", -- 7E00
         x"07",  x"03",  x"cb",  x"3e",  x"dc",  x"f6",  x"df",  x"1c", -- 7E08
         x"10",  x"f8",  x"c1",  x"d1",  x"e1",  x"3e",  x"f5",  x"3e", -- 7E10
         x"00",  x"32",  x"09",  x"03",  x"3e",  x"f5",  x"3e",  x"01", -- 7E18
         x"32",  x"08",  x"03",  x"f1",  x"c9",  x"7e",  x"fe",  x"23", -- 7E20
         x"20",  x"31",  x"cd",  x"bd",  x"c8",  x"30",  x"38",  x"23", -- 7E28
         x"e5",  x"e6",  x"03",  x"28",  x"12",  x"21",  x"07",  x"03", -- 7E30
         x"87",  x"fe",  x"04",  x"28",  x"12",  x"30",  x"16",  x"cb", -- 7E38
         x"4e",  x"cb",  x"ce",  x"20",  x"02",  x"c6",  x"08",  x"3c", -- 7E40
         x"32",  x"08",  x"03",  x"e1",  x"c3",  x"be",  x"c8",  x"cb", -- 7E48
         x"5e",  x"cb",  x"de",  x"18",  x"ee",  x"cb",  x"6e",  x"cb", -- 7E50
         x"ee",  x"18",  x"e8",  x"e5",  x"af",  x"18",  x"e8",  x"7e", -- 7E58
         x"fe",  x"23",  x"20",  x"30",  x"cd",  x"bd",  x"c8",  x"d2", -- 7E60
         x"48",  x"c3",  x"23",  x"e5",  x"e6",  x"03",  x"28",  x"12", -- 7E68
         x"21",  x"07",  x"03",  x"87",  x"fe",  x"04",  x"28",  x"10", -- 7E70
         x"38",  x"14",  x"cb",  x"66",  x"cb",  x"e6",  x"20",  x"02", -- 7E78
         x"c6",  x"08",  x"32",  x"09",  x"03",  x"e1",  x"18",  x"c4", -- 7E80
         x"cb",  x"56",  x"cb",  x"d6",  x"18",  x"f0",  x"cb",  x"46", -- 7E88
         x"cb",  x"c6",  x"18",  x"ea",  x"e5",  x"af",  x"18",  x"ea", -- 7E90
         x"c5",  x"cd",  x"2a",  x"d8",  x"e1",  x"23",  x"23",  x"23", -- 7E98
         x"23",  x"01",  x"61",  x"03",  x"c5",  x"18",  x"03",  x"cd", -- 7EA0
         x"d7",  x"de",  x"7e",  x"23",  x"fe",  x"22",  x"28",  x"16", -- 7EA8
         x"b7",  x"28",  x"1f",  x"f2",  x"a7",  x"de",  x"c5",  x"cd", -- 7EB0
         x"9a",  x"c7",  x"c1",  x"cd",  x"d7",  x"de",  x"1a",  x"13", -- 7EB8
         x"b7",  x"f2",  x"bb",  x"de",  x"18",  x"e4",  x"cd",  x"d7", -- 7EC0
         x"de",  x"7e",  x"23",  x"fe",  x"22",  x"28",  x"d8",  x"b7", -- 7EC8
         x"20",  x"f4",  x"3e",  x"20",  x"03",  x"18",  x"0c",  x"03", -- 7ED0
         x"02",  x"e5",  x"21",  x"56",  x"fc",  x"09",  x"e1",  x"d0", -- 7ED8
         x"e1",  x"3e",  x"2a",  x"cd",  x"d5",  x"dd",  x"af",  x"02", -- 7EE0
         x"e1",  x"77",  x"23",  x"e5",  x"cd",  x"f1",  x"c5",  x"d1", -- 7EE8
         x"23",  x"36",  x"00",  x"2b",  x"36",  x"20",  x"cd",  x"e4", -- 7EF0
         x"dd",  x"fe",  x"0a",  x"20",  x"05",  x"cd",  x"12",  x"df", -- 7EF8
         x"3c",  x"c9",  x"cd",  x"0f",  x"df",  x"c8",  x"cd",  x"27", -- 7F00
         x"df",  x"d8",  x"cd",  x"32",  x"df",  x"18",  x"e7",  x"fe", -- 7F08
         x"0d",  x"c0",  x"3e",  x"09",  x"cd",  x"d5",  x"dd",  x"23", -- 7F10
         x"7e",  x"b7",  x"20",  x"f6",  x"2b",  x"7e",  x"fe",  x"20", -- 7F18
         x"20",  x"02",  x"36",  x"00",  x"c3",  x"5e",  x"cb",  x"fe", -- 7F20
         x"03",  x"28",  x"02",  x"a7",  x"c9",  x"cd",  x"12",  x"df", -- 7F28
         x"37",  x"c9",  x"fe",  x"08",  x"28",  x"44",  x"fe",  x"09", -- 7F30
         x"28",  x"2a",  x"fe",  x"1f",  x"28",  x"47",  x"fe",  x"19", -- 7F38
         x"ca",  x"c5",  x"df",  x"fe",  x"18",  x"ca",  x"cf",  x"df", -- 7F40
         x"fe",  x"02",  x"ca",  x"db",  x"df",  x"fe",  x"1a",  x"28", -- 7F48
         x"48",  x"fe",  x"0b",  x"c8",  x"fe",  x"0a",  x"c8",  x"fe", -- 7F50
         x"01",  x"c8",  x"fe",  x"20",  x"30",  x"05",  x"3f",  x"cd", -- 7F58
         x"d5",  x"dd",  x"c9",  x"77",  x"cd",  x"d5",  x"dd",  x"23", -- 7F60
         x"7e",  x"b7",  x"c0",  x"11",  x"ab",  x"03",  x"cd",  x"89", -- 7F68
         x"c6",  x"28",  x"07",  x"36",  x"20",  x"23",  x"36",  x"00", -- 7F70
         x"18",  x"03",  x"cd",  x"a2",  x"c6",  x"2b",  x"7e",  x"b7", -- 7F78
         x"c0",  x"3e",  x"09",  x"18",  x"df",  x"e5",  x"23",  x"cd", -- 7F80
         x"f1",  x"c5",  x"cd",  x"a9",  x"c6",  x"d1",  x"af",  x"2b", -- 7F88
         x"46",  x"77",  x"cd",  x"a2",  x"c6",  x"78",  x"20",  x"f7", -- 7F90
         x"c9",  x"cd",  x"a9",  x"c6",  x"e5",  x"cd",  x"f1",  x"c5", -- 7F98
         x"11",  x"ab",  x"03",  x"cd",  x"89",  x"c6",  x"20",  x"0c", -- 7FA0
         x"cd",  x"a2",  x"c6",  x"cd",  x"a9",  x"c6",  x"cd",  x"a2", -- 7FA8
         x"c6",  x"2b",  x"36",  x"00",  x"d1",  x"44",  x"4d",  x"03", -- 7FB0
         x"7e",  x"02",  x"0b",  x"cd",  x"a2",  x"c6",  x"2b",  x"20", -- 7FB8
         x"f7",  x"23",  x"36",  x"20",  x"c9",  x"cd",  x"a2",  x"c6", -- 7FC0
         x"2b",  x"7e",  x"b7",  x"20",  x"f8",  x"18",  x"b2",  x"3e", -- 7FC8
         x"09",  x"cd",  x"d5",  x"dd",  x"23",  x"7e",  x"b7",  x"20", -- 7FD0
         x"f6",  x"18",  x"90",  x"cd",  x"c5",  x"df",  x"e5",  x"7e", -- 7FD8
         x"b7",  x"28",  x"05",  x"36",  x"20",  x"23",  x"18",  x"f7", -- 7FE0
         x"e1",  x"cd",  x"f1",  x"c5",  x"cd",  x"c5",  x"df",  x"23", -- 7FE8
         x"36",  x"00",  x"2b",  x"c9",  x"1e",  x"ff",  x"c3",  x"0e", -- 7FF0
         x"e0",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff"  -- 7FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
